problem "virtualhome-problem"
domain "virtualhome.cdl"

#!pragma planner_is_goal_serializable=False
#!pragma planner_is_goal_ordered=True
#!pragma planner_always_commit_skeleton=True

objects:
  light_1:item
  apple:item
  char:character

init:
  is_on[light_1] = True
  is_off[light_1] = False
  has_switch[light_1] = True
  sitting[char]=False
  close[char,light_1]=False
  holds_rh[char,apple]=False
  surfaces[light_1]=True
  grabbable[apple]=True
  inside[apple,light_1]=False
  inside[light_1,apple]=False
  on[apple,light_1]=False
  on[light_1,apple]=False

def dinner_prepared_for_two(coffe_maker_84: item):
  return is_on(coffe_maker_84)
  
behavior prepare_dinner_for_two(coffe_maker_84: item):
  goal:
    dinner_prepared_for_two(coffe_maker_84)
  body:
    achieve is_on(coffe_maker_84)

goal:
  on(apple,light_1)
