problem "kitchen-problem"
domain "kitchen_partial_ability.cdl"

#!pragma planner_is_goal_serializable=False
#!pragma planner_is_goal_ordered=True
#!pragma planner_always_commit_skeleton=True

objects:
#objects
  tomato_1:item
  tomato_2:item
  tomato_3:item
  tomato_4:item
  egg_5:item
  egg_6:item
  egg_7:item
  egg_8:item
  oil_9:item
  sugar_10:item
  pan_11:item
  salt_12:item
  bowl_13:item
  bowl_14:item
  bowl_15:item
  bowl_16:item
  knife_17:item
  fridge_18:item
  stove_19:item
  sink_20:item
  faucet_21:item
  spatula_22:item
  countertop_23:item
  water_24:item
  pepper_25:item
  bread_26:item
  onion_27:item
  bacon_28:item
  cheese_29:item
  bread_30:item
  bread_31:item
  bread_32:item
  pot_33:item
  noodles_34:item
  chicken_35:item
  garlic_36:item
  ginger_37:item
  vegetables_38:item
  oven_39:item
  plate_40:item
  plate_41:item
  plate_42:item
  plate_43:item
  cuttingboard_44:item
  beef_45:item
  potato_46:item
  shrimp_47:item

#object_end

init:
    #categories
    is_tomato[tomato_1]=True
    is_tomato[tomato_2]=True
    is_tomato[tomato_3]=True
    is_tomato[tomato_4]=True
    is_egg[egg_5]=True
    is_egg[egg_6]=True
    is_egg[egg_7]=True
    is_egg[egg_8]=True
    is_oil[oil_9]=True
    is_sugar[sugar_10]=True
    is_pan[pan_11]=True
    is_salt[salt_12]=True
    is_bowl[bowl_13]=True
    is_bowl[bowl_14]=True
    is_bowl[bowl_15]=True
    is_bowl[bowl_16]=True
    is_plate[plate_40]=True
    is_plate[plate_41]=True
    is_plate[plate_42]=True
    is_plate[plate_43]=True
    is_knife[knife_17]=True
    is_fridge[fridge_18]=True
    is_stove[stove_19]=True
    is_sink[sink_20]=True
    is_faucet[faucet_21]=True
    is_spatula[spatula_22]=True
    is_countertop[countertop_23]=True
    is_water[water_24]=True
    is_pepper[pepper_25]=True
    is_bread[bread_26]=True
    is_onion[onion_27]=True
    is_bacon[bacon_28]=True
    is_cheese[cheese_29]=True
    is_bread[bread_30]=True
    is_bread[bread_31]=True
    is_bread[bread_32]=True
    is_pot[pot_33]=True
    is_noodles[noodles_34]=True
    is_chicken[chicken_35]=True
    is_garlic[garlic_36]=True
    is_ginger[ginger_37]=True
    is_vegetables[vegetables_38]=True
    is_oven[oven_39]=True
    is_cuttingboard[cuttingboard_44]=True
    is_beef[beef_45]=True
    is_potato[potato_46]=True
    is_shrimp[shrimp_47]=True
    #categories_end

    #states
    is_off[stove_19]=True
    is_on[stove_19]=False
    is_off[faucet_21]=True
    is_on[faucet_21]=False
    is_off[oven_39]=True
    is_on[oven_39]=False
    open[fridge_18]=False
    closed[fridge_18]=True
    open[oven_39]=False
    closed[oven_39]=True
    dirty[pan_11]=False
    clean[pan_11]=True
    dirty[pot_33]=False
    clean[pot_33]=True
    dirty[bowl_13]=False
    clean[bowl_13]=True
    dirty[bowl_14]=False
    clean[bowl_14]=True
    dirty[bowl_15]=False
    clean[bowl_15]=True
    dirty[bowl_16]=False
    clean[bowl_16]=True
    dirty[plate_40]=False
    clean[plate_40]=True
    dirty[plate_41]=False
    clean[plate_41]=True
    dirty[plate_42]=False
    clean[plate_42]=True
    dirty[plate_43]=False
    clean[plate_43]=True
    dirty[tomato_1]=True
    clean[tomato_1]=False
    dirty[tomato_2]=True
    clean[tomato_2]=False
    dirty[tomato_3]=True
    clean[tomato_3]=False
    dirty[tomato_4]=True
    clean[tomato_4]=False
    sliced[tomato_1]=False
    sliced[tomato_2]=False
    sliced[tomato_3]=False
    sliced[tomato_4]=False
    dirty[onion_27]=True
    clean[onion_27]=False
    dirty[vegetables_38]=True
    clean[vegetables_38]=False
    peeled[onion_27]=False
    sliced[onion_27]=False
    peeled[egg_5]=False
    peeled[egg_6]=False
    peeled[egg_7]=False
    peeled[egg_8]=False
    peeled[tomato_1]=False
    peeled[tomato_2]=False
    peeled[tomato_3]=False
    peeled[tomato_4]=False
    mixed[bowl_13]=False
    mixed[bowl_14]=False
    mixed[bowl_15]=False
    mixed[bowl_16]=False
    mixed[pan_11]=False
    mixed[pot_33]=False
    waterfull[sink_20]=False
    waterfull[pan_11]=False
    waterfull[pot_33]=False
    waterfull[bowl_13]=False
    waterfull[bowl_14]=False
    waterfull[bowl_15]=False
    waterfull[bowl_16]=False
    #states_end

    #properties
    surfaces[countertop_23]=True
    surfaces[stove_19]=True
    surfaces[cuttingboard_44]=True
    grabbable[tomato_1]=True
    grabbable[tomato_2]=True
    grabbable[tomato_3]=True
    grabbable[tomato_4]=True
    grabbable[egg_5]=True
    grabbable[egg_6]=True
    grabbable[egg_7]=True
    grabbable[egg_8]=True
    grabbable[oil_9]=True
    grabbable[sugar_10]=True
    grabbable[pan_11]=True
    grabbable[salt_12]=True
    grabbable[bowl_13]=True
    grabbable[bowl_14]=True
    grabbable[bowl_15]=True
    grabbable[bowl_16]=True
    grabbable[knife_17]=True
    grabbable[spatula_22]=True
    grabbable[pepper_25]=True
    grabbable[bread_26]=True
    grabbable[onion_27]=True
    grabbable[bacon_28]=True
    grabbable[cheese_29]=True
    grabbable[bread_30]=True
    grabbable[bread_31]=True
    grabbable[bread_32]=True
    grabbable[pot_33]=True
    grabbable[noodles_34]=True
    grabbable[chicken_35]=True
    grabbable[garlic_36]=True
    grabbable[ginger_37]=True
    grabbable[vegetables_38]=True
    grabbable[plate_40]=True
    grabbable[plate_41]=True
    grabbable[plate_42]=True
    grabbable[plate_43]=True
    grabbable[cuttingboard_44]=True
    grabbable[beef_45]=True
    grabbable[potato_46]=True
    grabbable[shrimp_47]=True
    cuttable[tomato_1]=True
    cuttable[tomato_2]=True
    cuttable[tomato_3]=True
    cuttable[tomato_4]=True
    cuttable[onion_27]=True
    cuttable[cheese_29]=True
    cuttable[bacon_28]=True
    cuttable[bread_26]=True
    cuttable[bread_30]=True
    cuttable[bread_31]=True
    cuttable[bread_32]=True
    cuttable[noodles_34]=True
    cuttable[chicken_35]=True
    cuttable[garlic_36]=True
    cuttable[ginger_37]=True
    cuttable[vegetables_38]=True
    cuttable[beef_45]=True
    cuttable[potato_46]=True
    cuttable[shrimp_47]=True
    containers[fridge_18]=True
    containers[bowl_13]=True
    containers[bowl_14]=True
    containers[bowl_15]=True
    containers[bowl_16]=True
    containers[plate_40]=True
    containers[plate_41]=True
    containers[plate_42]=True
    containers[plate_43]=True
    containers[pan_11]=True
    containers[pot_33]=True
    containers[sink_20]=True
    containers[oven_39]=True
    peelable[tomato_1]=True
    peelable[tomato_2]=True
    peelable[tomato_3]=True
    peelable[tomato_4]=True
    peelable[potato_46]=True
    peelable[shrimp_47]=True
    can_open[fridge_18]=True
    can_open[oven_39]=True
    has_switch[stove_19]=True
    has_switch[faucet_21]=True
    has_switch[oven_39]=True
    eatable[tomato_1]=True
    eatable[tomato_2]=True
    eatable[tomato_3]=True
    eatable[tomato_4]=True
    eatable[egg_5]=True
    eatable[egg_6]=True
    eatable[egg_7]=True
    eatable[egg_8]=True
    eatable[oil_9]=True
    eatable[sugar_10]=True
    eatable[salt_12]=True
    eatable[pepper_25]=True
    eatable[bread_26]=True
    eatable[onion_27]=True
    eatable[bacon_28]=True
    eatable[cheese_29]=True
    eatable[bread_30]=True
    eatable[bread_31]=True
    eatable[bread_32]=True
    eatable[noodles_34]=True
    eatable[chicken_35]=True
    eatable[garlic_36]=True
    eatable[ginger_37]=True
    eatable[vegetables_38]=True
    eatable[beef_45]=True
    eatable[potato_46]=True
    eatable[shrimp_47]=True
    cookaware[pan_11]=True
    cookaware[pot_33]=True
    cookaware[oven_39]=True
    storable[countertop_23]=True
    pourable[pepper_25]=True
    pourable[salt_12]=True
    #properties_end

    #relations
    inside[tomato_1,fridge_18]=True
    inside[tomato_2,fridge_18]=True
    inside[tomato_3,fridge_18]=True
    inside[tomato_4,fridge_18]=True
    close[tomato_1,fridge_18]=True
    close[tomato_2,fridge_18]=True
    close[tomato_3,fridge_18]=True
    close[tomato_4,fridge_18]=True
    close[fridge_18,tomato_1]=True
    close[fridge_18,tomato_2]=True
    close[fridge_18,tomato_3]=True
    close[fridge_18,tomato_4]=True
    inside[egg_5,fridge_18]=True
    inside[egg_6,fridge_18]=True
    inside[egg_7,fridge_18]=True
    inside[egg_8,fridge_18]=True
    close[egg_5,fridge_18]=True
    close[egg_6,fridge_18]=True
    close[egg_7,fridge_18]=True
    close[egg_8,fridge_18]=True
    close[fridge_18,egg_5]=True
    close[fridge_18,egg_6]=True
    close[fridge_18,egg_7]=True
    close[fridge_18,egg_8]=True
    inside[bread_26,fridge_18]=True
    close[bread_26,fridge_18]=True
    close[fridge_18,bread_26]=True
    inside[bread_30,fridge_18]=True
    close[bread_30,fridge_18]=True
    close[fridge_18,bread_30]=True
    inside[bread_31,fridge_18]=True
    close[bread_31,fridge_18]=True
    close[fridge_18,bread_31]=True
    inside[bread_32,fridge_18]=True
    close[bread_32,fridge_18]=True
    close[fridge_18,bread_32]=True
    inside[onion_27,fridge_18]=True
    close[onion_27,fridge_18]=True
    close[fridge_18,onion_27]=True
    inside[bacon_28,fridge_18]=True
    close[bacon_28,fridge_18]=True
    close[fridge_18,bacon_28]=True
    inside[cheese_29,fridge_18]=True
    close[cheese_29,fridge_18]=True
    close[fridge_18,cheese_29]=True
    inside[noodles_34,fridge_18]=True
    close[noodles_34,fridge_18]=True
    close[fridge_18,noodles_34]=True
    on[pan_11,countertop_23]=True
    close[pan_11,countertop_23]=True
    close[countertop_23,pan_11]=True
    on[pot_33,countertop_23]=True
    close[pot_33,countertop_23]=True
    close[countertop_23,pot_33]=True
    on[faucet_21,sink_20]=True
    close[faucet_21,sink_20]=True
    close[sink_20,faucet_21]=True
    on[bowl_13,countertop_23]=True
    close[bowl_13,countertop_23]=True
    close[countertop_23,bowl_13]=True
    on[bowl_14,countertop_23]=True
    close[bowl_14,countertop_23]=True
    close[countertop_23,bowl_14]=True
    on[bowl_15,countertop_23]=True
    close[bowl_15,countertop_23]=True
    close[countertop_23,bowl_15]=True
    on[bowl_16,countertop_23]=True
    close[bowl_16,countertop_23]=True
    close[countertop_23,bowl_16]=True
    on[plate_40,countertop_23]=True
    close[plate_40,countertop_23]=True
    close[countertop_23,plate_40]=True
    on[plate_41,countertop_23]=True
    close[plate_41,countertop_23]=True
    close[countertop_23,plate_41]=True
    on[plate_42,countertop_23]=True
    close[plate_42,countertop_23]=True
    close[countertop_23,plate_42]=True
    on[plate_43,countertop_23]=True
    close[plate_43,countertop_23]=True
    close[countertop_23,plate_43]=True
    inside[spatula_22,pan_11]=True
    close[spatula_22,pan_11]=True
    close[pan_11,spatula_22]=True
    on[knife_17,countertop_23]=True
    close[knife_17,countertop_23]=True
    close[countertop_23,knife_17]=True
    on[oil_9,countertop_23]=True
    close[oil_9,countertop_23]=True
    close[countertop_23,oil_9]=True
    on[sugar_10,countertop_23]=True
    close[sugar_10,countertop_23]=True
    close[countertop_23,sugar_10]=True
    on[salt_12,countertop_23]=True
    close[salt_12,countertop_23]=True
    close[countertop_23,salt_12]=True
    on[pepper_25,countertop_23]=True
    close[pepper_25,countertop_23]=True
    close[countertop_23,pepper_25]=True
    on[garlic_36,countertop_23]=True
    close[garlic_36,countertop_23]=True
    close[countertop_23,garlic_36]=True
    on[ginger_37,countertop_23]=True
    close[ginger_37,countertop_23]=True
    close[countertop_23,ginger_37]=True
    inside[vegetables_38,fridge_18]=True
    close[vegetables_38,fridge_18]=True
    close[fridge_18,vegetables_38]=True
    inside[chicken_35,fridge_18]=True
    close[chicken_35,fridge_18]=True
    close[fridge_18,chicken_35]=True
    on[oven_39,countertop_23]=True
    close[oven_39,countertop_23]=True
    close[countertop_23,oven_39]=True
    on[cuttingboard_44,countertop_23]=True
    close[cuttingboard_44,countertop_23]=True
    close[countertop_23,cuttingboard_44]=True
    inside[beef_45,fridge_18]=True
    close[beef_45,fridge_18]=True
    close[fridge_18,beef_45]=True
    inside[potato_46,fridge_18]=True
    close[potato_46,fridge_18]=True
    close[fridge_18,potato_46]=True
    inside[shrimp_47,fridge_18]=True
    close[shrimp_47,fridge_18]=True
    close[fridge_18,shrimp_47]=True
    #relations_end

    #id
    id[tomato_1]=1
    id[tomato_2]=2
    id[tomato_3]=3
    id[tomato_4]=4
    id[egg_5]=5
    id[egg_6]=6
    id[egg_7]=7
    id[egg_8]=8
    id[oil_9]=9
    id[sugar_10]=10
    id[pan_11]=11
    id[salt_12]=12
    id[bowl_13]=13
    id[bowl_14]=14
    id[bowl_15]=15
    id[bowl_16]=16
    id[knife_17]=17
    id[fridge_18]=18
    id[stove_19]=19
    id[sink_20]=20
    id[faucet_21]=21
    id[spatula_22]=22
    id[countertop_23]=23
    id[water_24]=24
    id[pepper_25]=25
    id[bread_26]=26
    id[onion_27]=27
    id[bacon_28]=28
    id[cheese_29]=29
    id[bread_30]=30
    id[bread_31]=31
    id[bread_32]=32
    id[pot_33]=33
    id[noodles_34]=34
    id[chicken_35]=35
    id[garlic_36]=36
    id[ginger_37]=37
    id[vegetables_38]=38
    id[oven_39]=39
    id[plate_40]=40
    id[plate_41]=41
    id[plate_42]=42
    id[plate_43]=43
    id[cuttingboard_44]=44
    id[beef_45]=45
    id[potato_46]=46
    id[shrimp_47]=47
    #id_end

#exploration
    known[fridge_18]=True
    known[stove_19]=True
    known[sink_20]=True
    known[faucet_21]=True
    known[countertop_23]=True
    known[oven_39]=True
    #exploration_end

