problem "agent-problem"
domain "virtualhome_partial.cdl"

objects:
  cup_a: item
  cup_b: item

init:
  is_cup[cup_a] = True
  is_cup[cup_b] = True
  grabbable[cup_a] = False
  grabbable[cup_b] = True
  has_a_free_hand[char] = True

behavior get_a_cup():
  body:
    bind cup: item where:
      is_cup(cup)
    achieve inhand(cup)

behavior __goal__():
  body:
    get_a_cup()
      
  