
behavior heat_in_microwave(plate:item, microwave:item):
    body:
        achieve_once inside(plate, microwave)
        # Place the plate inside the microwave
        achieve_once closed(microwave)
        # Close the microwave
        achieve_once is_on(microwave)
        # Turn on the microwave

behavior __goal__():
    body:
        bind plate: item where:
            is_plate(plate) and on(food_pizza_2065, plate) and on(food_hamburger_2057, plate)
        # Select the plate with both pizza and hamburger on it

        bind microwave: item where:
            is_microwave(microwave)
        # Select a microwave

        heat_in_microwave(plate, microwave)
        # Heat the plate with pizza and hamburger in the microwave
