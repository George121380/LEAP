problem "agent-problem"
domain "virtualhome_partial.cdl"

objects:
  cup_a: item
  cup_b: item
  fridge: item

init:
  is_cup[cup_a] = True
  is_cup[cup_b] = True
  is_fridge[fridge] = True
  grabbable[cup_a] = True
  grabbable[cup_b] = True
  containers[fridge] = True
  has_a_free_hand[char] = True
  size[cup_a] = 10
  size[cup_b] = 5
  size[fridge] = 8
  close_char[char,fridge] = False

behavior __goal__():
  body:
    bind f: item where:
      is_fridge(f)
    bind c: item where:
      is_cup(c)
    achieve inside(c,f)
      
  