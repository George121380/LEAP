 
behavior cook_chicken(chicken:item, stove:item):
    body:
        achieve on(chicken, stove)
        achieve is_on(stove)

behavior cook_pasta(pasta:item, pot:item, stove:item):
    body:
        achieve inside(pasta, pot)
        achieve on(pot, stove)
        achieve is_on(stove)

behavior __goal__():
    body:
        bind stove: item where:
            is_stove(stove)
        # Select the stove

        bind chicken: item where:
            is_food_chicken(chicken)
        # Select the chicken

        bind pot: item where:
            is_pot(pot)
        # Select the pot
        
        bind pasta: item where:
            is_dry_pasta(pasta)
        # Select the pasta

        cook_chicken(chicken, stove)
        cook_pasta(pasta, pot, stove)
