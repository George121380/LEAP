 
behavior find_book_and_put_on_table(book:item, table:item):
    body:
        achieve inside(book, table)
        # Ensure the book is placed on the table

behavior turn_on_light(light:item):
    body:
        achieve is_on(light)
        # Turn on the light

behavior __goal__():
    body:
        bind home_office: item where:
            is_home_office(home_office)
        # Select the home office

        bind book: item where:
            is_book(book)
        # Select a book

        bind table: item where:
            is_table(table) and inside(table, home_office)
        # Select a table inside the home office

        bind light: item where:
            is_light(light) and inside(light, home_office)
        # Select a light inside the home office

        find_book_and_put_on_table(book, table)
        turn_on_light(light)
