problem "virtualhome-problem"
domain "virtualhome.cdl"

#!pragma planner_is_goal_serializable=False
#!pragma planner_is_goal_ordered=True
#!pragma planner_always_commit_skeleton=True

objects:
  light:item
  char:character
  apple:item

init:
  is_on[light] = True
  is_off[light] = False
  sitting[char]=False
  lying[char]=False
  close[char,light]=False
  holds_rh[char,apple]=False
  surfaces[light]=True
  grabbable[apple]=True



goal:
  on(apple,light)
