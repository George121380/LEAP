typedef Object: object

feature is_object(x: Object) -> bool
feature is_container(x: Object) -> bool
feature can_contain(x: Object, y: Object) -> bool

feature contained_in_something(x: Object) -> bool # x is contained in something
feature containing(c: Object, x: Object) -> bool # x is contained in c

controller put_into(x: Object, y: Object)

behavior put_object_into_container(x: Object):
    goal: contained_in_something(x)
    body:
        bind c: Object where: (
            is_container(c) and
            can_contain(c, x) and
            not (exists y: Object: containing(c, y))
        )
        put_into(x, c)
    eff:
        contained_in_something[x] = True
        containing[c, x] = True