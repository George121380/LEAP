domain "virtualhome"

typedef item: object
typedef character: object

# Features without return type annotations are assumed to be returning boolean values.

#state
feature is_on(x: item)
feature is_off(x: item)
feature plugged(x: item)
feature unplugged(x: item)
feature open(x: item)
feature closed(x: item)
feature dirty(x: item)
feature clean(x: item)
feature sitting(x: character)
feature lying(x: character)

#add state
feature is_room(x: item)

#relationship
feature on(x: item, y: item)
feature on_char(x: character, y: item)
feature inside(x: item, y: item)
feature inside_char(x: character, y: item)

feature between(door: item, room: item)
feature close_item(x: item, y: item)
feature close(x: character, y: item)
feature facing_item(x: item, y: item)
feature facing(x: character, y: item)
feature holds_rh(x: character, y: item)
feature holds_lh(x: character, y: item)

#Properties 
feature surfaces(x: item)
feature grabbable(x: item)
feature sittable(x: item)
feature lieable(x: item)
feature hangable(x: item)
feature drinkable(x: item)
feature eatable(x: item)
feature recipient(x: item)
feature cuttable(x: item)
feature pourable(x: item)
feature can_open(x: item)
feature has_switch(x: item)
feature readable(x: item)
feature lookable(x: item)
feature containers(x: item)
feature clothes(x: item)
feature person(x: item)
feature body_part(x: item)
feature cover_object(x: item)
feature has_plug(x: item)
feature has_paper(x: item)
feature movable(x: item)
feature cream(x: item)


object_constant char:character

#controllers
controller walk_executor(x: item)
controller switchoff_executor(x: item)
controller switchon_executor(x: item)
controller put_executor(x: item, y: item)
controller grab_executor(x: item)
controller standup_executor(x: character)
controller wash_executor(x: item)
controller sit_executor(x: character)
controller open_executor(x: item)
controller close_executor(x: item)
controller pour_executor(x: item, y: item)
controller plugin_executor(x: item)
controller plugout_executor(x: item)


def inhand(inhand_obj:item):
  return holds_rh(char, inhand_obj) or holds_lh(char, inhand_obj)

def standing(char: character):
  return not sitting(char) and not lying(char)

def has_a_free_hand():
  symbol l=exists item1: item : holds_lh(char, item1)
  symbol r=exists item2: item : holds_rh(char, item2)
  return not l or not r



behavior put(inhand_obj: item, obj: item):
  body:
    assert surfaces(obj)
    achieve inhand(inhand_obj)
    achieve close(char, obj)
    put_executor(inhand_obj, obj)
  eff:
    holds_rh[char, inhand_obj] = False
    holds_lh[char, inhand_obj] = False
    on[inhand_obj, obj] = True
    close_item[inhand_obj, obj] = True
    close_item[obj, inhand_obj] = True
    foreach inter:item:
      if close_item(inter, obj):
        close_item[inter, inhand_obj] = True
        close_item[inhand_obj, inter] = True

behavior empty_a_hand():
  goal: has_a_free_hand()
  body:
    assert not has_a_free_hand()
    bind surf:item where:
      surfaces(surf)
    bind give_up_obj:item where:
      inhand(give_up_obj)
    put(give_up_obj, surf)

behavior stand():
  goal: standing(char)
  body:
    assert sitting(char) or lying(char)
    standup_executor(char)
  eff:
    sitting[char] = False
    lying[char] = False

behavior sit(obj: item):
  goal: sitting(char)
  body:
    assert sittable(obj)
    assert not sitting(char)
    achieve close(char, obj)
    sit_executor(char)
  eff:
    sitting[char] = True
    on_char[char, obj] = True

def obj_inside_or_on(obj1: item, obj2: item):
  return inside(obj1, obj2) or on(obj2, obj1)

behavior walk(obj: item):
  goal: close(char, obj)
  body:
    achieve standing(char)
    walk_executor(obj)
  eff:
    foreach icf:item:
      close[char, icf]= False
      facing[char, icf]= False
      inside_char[char,icf]= False
      if obj_inside_or_on(obj, icf):
        close[char, icf] = True
    close[char,obj] = True

behavior switch_off(obj: item):
  goal: is_off(obj)
  body:
    assert has_switch(obj)
    assert is_on(obj)
    achieve has_a_free_hand()
    achieve close(char, obj)
    switchoff_executor(obj)
  eff:
    is_off[obj] = True
    is_on[obj] = False

behavior switch_on(obj: item):
  goal: is_on(obj)
  body:
    assert has_switch(obj)
    assert is_off(obj)
    achieve has_a_free_hand()
    achieve close(char, obj)
    switchon_executor(obj)
  eff:
    is_off[obj] = False
    is_on[obj] = True

behavior put_close(inhand_obj: item, obj: item):
  goal: close_item(inhand_obj, obj)
  body:
    put(inhand_obj, obj)

behavior put_on(inhand_obj: item, obj: item):
  goal: on(inhand_obj, obj)
  body:
    put(inhand_obj, obj)

behavior grab(obj: item):
  goal: inhand(obj)
  body:
    assert grabbable(obj)
    achieve has_a_free_hand()
    foreach obj2:item:
      if inside(obj,obj2):
        if not is_room(obj2):
          assert can_open(obj2)
          achieve open(obj2)
    achieve close(char, obj)
    grab_executor(obj)
  eff:
    holds_rh[char,obj]=True

behavior wash(obj: item):
  goal: clean(obj)
  body:
    achieve has_a_free_hand()
    achieve close(char, obj)
    wash_executor(obj)
  eff:
    dirty[obj] = False
    clean[obj] = True

behavior open(obj: item):
  goal: open(obj)
  body:
    assert can_open(obj)
    assert closed(obj)
    achieve has_a_free_hand()
    achieve close(char, obj)
    open_executor(obj)
  eff:
    open[obj] = True
    closed[obj] = False

behavior close(obj: item):
  goal: closed(obj)
  body:
    assert can_open(obj)
    assert open(obj)
    achieve has_a_free_hand()
    achieve close(char, obj)
    close_executor(obj)
  eff:
    open[obj] = False
    closed[obj] = True

behavior pour(obj: item, target: item):
  goal: inside(obj, target)
  body:
    assert pourable(obj) or drinkable(obj)
    assert recipient(target)
    achieve inhand(obj)
    achieve close(char, target)
    pour_executor(obj, target)
  eff:
    inside[obj, target] = True

behavior plugin(object:item):
  goal: plugged(object)
  body:
    assert has_plug(object)
    assert unplugged(object)
    achieve has_a_free_hand()
    achieve close(char, object)
    plugin_executor(object)
  eff:
    plugged[object] = True
    unplugged[object] = False
  
behavior plugout(object:item):
  goal: unplugged(object)
  body:
    assert has_plug(object)
    assert plugged(object)
    achieve has_a_free_hand()
    achieve close(char, object)
    plugout_executor(object)
  eff:
    plugged[object] = False
    unplugged[object] = True