domain "virtualhome_partial"

typedef item: object
typedef character: object
typedef id: int64
# Features without return type annotations are assumed to be returning boolean values.

#state
feature is_on(x: item)
feature is_off(x: item)
feature plugged(x: item)
feature unplugged(x: item)
feature open(x: item)
feature closed(x: item)
feature dirty(x: item)
feature clean(x: item)
feature sitting(x: character)
feature lying(x: character)
feature standing(x: character)
feature cut(x:item)
feature sleeping(x: character)
feature inhand(x: item)
feature visited(x: item)
feature has_water(x: item)
feature used(x: item)
feature has_a_free_hand(x: character)

#relationship
feature on(x: item, y: item)
feature inside(x: item, y: item)
feature between(door: item, room: item)
feature close(x: item, y: item)
feature facing(x: item, y: item)
feature close_char(x: character, y: item)
feature facing_char(x: character, y: item)
feature inside_char(x: character, y: item)
feature on_char(x: character, y: item)
feature on_body(x:item, y: character)
feature holds_rh(x: character, y: item)
feature holds_lh(x: character, y: item)

#Properties
feature surfaces(x: item)
feature grabbable(x: item)
feature sittable(x: item)
feature lieable(x: item)
feature hangable(x: item)
feature drinkable(x: item)
feature eatable(x: item)
feature recipient(x: item)
feature cuttable(x: item)
feature pourable(x: item)
feature can_open(x: item)
feature has_switch(x: item)
feature readable(x: item)
feature lookable(x: item)
feature containers(x: item)
feature person(x: item)
feature body_part(x: item)
feature cover_object(x: item)
feature has_plug(x: item)
feature has_paper(x: item)
feature movable(x: item)
feature cream(x: item)
feature is_clothes(x: item)
feature is_food(x: item)
feature has_size(x: item)

object_constant char:character

feature id(x:item) -> int64
feature size(x:item) -> int64

#exploration
feature unknown(x: item)

#category
feature is_carrot(x:item)
feature is_candle(x:item)
feature is_coin(x:item)
feature is_dishwashingliquid(x:item)
feature is_balanceball(x:item)
feature is_cleaning_bottle(x:item)
feature is_bellpepper(x:item)
feature is_blow_dryer(x:item)
feature is_coffee_table(x:item)
feature is_food_bacon(x:item)
feature is_cpu_case(x:item)
feature is_crayon(x:item)
feature is_food_carrot(x:item)
feature is_ground_coffee(x:item)
feature is_bread(x:item)
feature is_drinking_glass(x:item)
feature is_scissors(x:item)
feature is_thread(x:item)
feature is_sauce_pan(x:item)
feature is_mincedmeat(x:item)
feature is_food_pizza(x:item)
feature is_oil(x:item)
feature is_walltv(x:item)
feature is_dirt(x:item)
feature is_cpu_table(x:item)
feature is_food_fruit(x:item)
feature is_music_stand(x:item)
feature is_living_room(x:item)
feature is_lamp(x:item)
feature is_clock(x:item)
feature is_bathroom_counter(x:item)
feature is_chefknife(x:item)
feature is_man(x:item)
feature is_tea(x:item)
feature is_bag(x:item)
feature is_salmon(x:item)
feature is_food_salt(x:item)
feature is_globe(x:item)
feature is_picture(x:item)
feature is_food_cereal(x:item)
feature is_duster(x:item)
feature is_juice(x:item)
feature is_clothes_socks(x:item)
feature is_room(x:item)
feature is_wine_glass(x:item)
feature is_chinesefood(x:item)
feature is_broom(x:item)
feature is_kettle(x:item)
feature is_light_bulb(x:item)
feature is_bucket(x:item)
feature is_sink(x:item)
feature is_faucet(x:item)
feature is_milkshake(x:item)
feature is_mouthwash(x:item)
feature is_comb(x:item)
feature is_mail(x:item)
feature is_glasses(x:item)
feature is_envelope(x:item)
feature is_tvstand(x:item)
feature is_newspaper(x:item)
feature is_washing_sponge(x:item)
feature is_printer(x:item)
feature is_purse(x:item)
feature is_toaster(x:item)
feature is_toy(x:item)
feature is_dvd_player(x:item)
feature is_rug(x:item)
feature is_bottle_water(x:item)
feature is_tooth_paste(x:item)
feature is_clothes_pile(x:item)
feature is_clothes_pants(x:item)
feature is_mat(x:item)
feature is_coffee_filter(x:item)
feature is_knifeblock(x:item)
feature is_toiletpaper(x:item)
feature is_curtain(x:item)
feature is_food_sugar(x:item)
feature is_kitchen_counter(x:item)
feature is_plate(x:item)
feature is_measuring_cup(x:item)
feature is_fax_machine(x:item)
feature is_creditcard(x:item)
feature is_closet(x:item)
feature is_kitchen_cabinets(x:item)
feature is_orchid(x:item)
feature is_cloth_napkin(x:item)
feature is_fryingpan(x:item)
feature is_bathtub(x:item)
feature is_toothpaste(x:item)
feature is_electric_shaver(x:item)
feature is_pear(x:item)
feature is_stove(x:item)
feature is_mop(x:item)
feature is_water_glass(x:item)
feature is_ice(x:item)
feature is_cat(x:item)
feature is_centerpiece(x:item)
feature is_face_cream(x:item)
feature is_food_potato(x:item)
feature is_food_oatmeal(x:item)
feature is_dishrack(x:item)
feature is_console(x:item)
feature is_hairdryer(x:item)
feature is_nightstand(x:item)
feature is_facial_cleanser(x:item)
feature is_detergent(x:item)
feature is_jelly(x:item)
feature is_chair(x:item)
feature is_sheets(x:item)
feature is_dustpan(x:item)
feature is_tablelamp(x:item)
feature is_novel(x:item)
feature is_mug(x:item)
feature is_entrance_hall(x:item)
feature is_phone(x:item)
feature is_cutting_board(x:item)
feature is_coffeetable(x:item)
feature is_cd(x:item)
feature is_lighter(x:item)
feature is_microwave(x:item)
feature is_dishwasher(x:item)
feature is_hairproduct(x:item)
feature is_food_turkey(x:item)
feature is_stamp(x:item)
feature is_wall_phone(x:item)
feature is_bookmark(x:item)
feature is_colander(x:item)
feature is_carpet(x:item)
feature is_glass(x:item)
feature is_ceilinglamp(x:item)
feature is_scrabble(x:item)
feature is_food_hamburger(x:item)
feature is_clothes_scarf(x:item)
feature is_fly(x:item)
feature is_clothes_jacket(x:item)
feature is_cucumber(x:item)
feature is_cookingpot(x:item)
feature is_document(x:item)
feature is_food_lime(x:item)
feature is_laser_pointer(x:item)
feature is_food_butter(x:item)
feature is_cards(x:item)
feature is_tray(x:item)
feature is_fork(x:item)
feature is_face_soap(x:item)
feature is_notes(x:item)
feature is_dog(x:item)
feature is_potato(x:item)
feature is_food_ice_cream(x:item)
feature is_teddybear(x:item)
feature is_oventray(x:item)
feature is_instrument_violin(x:item)
feature is_kitchen_cabinet(x:item)
feature is_oven_mitts(x:item)
feature is_nail_polish(x:item)
feature is_pot(x:item)
feature is_address_book(x:item)
feature is_wine(x:item)
feature is_food_donut(x:item)
feature is_table_cloth(x:item)
feature is_cd_player(x:item)
feature is_cutlery_knife(x:item)
feature is_clothes_shirt(x:item)
feature is_slippers(x:item)
feature is_cooking_pot(x:item)
feature is_mousemat(x:item)
feature is_television(x:item)
feature is_ironing_board(x:item)
feature is_cpuscreen(x:item)
feature is_shower(x:item)
feature is_coffee(x:item)
feature is_fridge(x:item)
feature is_shoe_shine_kit(x:item)
feature is_magazine(x:item)
feature is_food_food(x:item)
feature is_light(x:item)
feature is_book(x:item)
feature is_painting(x:item)
feature is_towel_rack(x:item)
feature is_food_noodles(x:item)
feature is_food_rice(x:item)
feature is_coffe_maker(x:item)
feature is_ceilingfan(x:item)
feature is_sportsball(x:item)
feature is_clothes_skirt(x:item)
feature is_light_switch(x:item)
feature is_window(x:item)
feature is_walllamp(x:item)
feature is_shredder(x:item)
feature is_filing_cabinet(x:item)
feature is_keys(x:item)
feature is_mirror(x:item)
feature is_chef_knife(x:item)
feature is_laundry_detergent(x:item)
feature is_salt_crackers(x:item)
feature is_iron(x:item)
feature is_drying_rack(x:item)
feature is_face(x:item)
feature is_clothes_gloves(x:item)
feature is_banana(x:item)
feature is_tomato(x:item)
feature is_dough(x:item)
feature is_orange(x:item)
feature is_bowl(x:item)
feature is_printing_paper(x:item)
feature is_sponge(x:item)
feature is_longboard(x:item)
feature is_coffee_cup(x:item)
feature is_check(x:item)
feature is_video_game_console(x:item)
feature is_drawing(x:item)
feature is_controller(x:item)
feature is_beer(x:item)
feature is_photoframe(x:item)
feature is_floor_lamp(x:item)
feature is_watermelon(x:item)
feature is_bathroom(x:item)
feature is_shoe_rack(x:item)
feature is_mouse(x:item)
feature is_deck_of_cards(x:item)
feature is_shaving_cream(x:item)
feature is_mechanical_pencil(x:item)
feature is_milk(x:item)
feature is_bathroom_cabinet(x:item)
feature is_waterglass(x:item)
feature is_toilet(x:item)
feature is_needle(x:item)
feature is_tape(x:item)
feature is_pc(x:item)
feature is_apple(x:item)
feature is_shampoo(x:item)
feature is_freezer(x:item)
feature is_trashcan(x:item)
feature is_alcohol(x:item)
feature is_pasta(x:item)
feature is_basket_for_clothes(x:item)
feature is_condiment_shaker(x:item)
feature is_toilet_paper(x:item)
feature is_barsoap(x:item)
feature is_food_jam(x:item)
feature is_napkin(x:item)
feature is_food_dessert(x:item)
feature is_brush(x:item)
feature is_mousepad(x:item)
feature is_feet_both(x:item)
feature is_chicken(x:item)
feature is_hairbrush(x:item)
feature is_boardgame(x:item)
feature is_cleaning_solution(x:item)
feature is_sofa(x:item)
feature is_wallpictureframe(x:item)
feature is_button(x:item)
feature is_coatrack(x:item)
feature is_pillow(x:item)
feature is_spoon(x:item)
feature is_bed(x:item)
feature is_blanket(x:item)
feature is_lightswitch(x:item)
feature is_radio(x:item)
feature is_stereo(x:item)
feature is_cutlets(x:item)
feature is_whippedcream(x:item)
feature is_water(x:item)
feature is_headset(x:item)
feature is_bookshelf(x:item)
feature is_clothes_hat(x:item)
feature is_cabinet(x:item)
feature is_hanger(x:item)
feature is_food_egg(x:item)
feature is_standingmirror(x:item)
feature is_knife(x:item)
feature is_stovefan(x:item)
feature is_food_kiwi(x:item)
feature is_vase(x:item)
feature is_wallshelf(x:item)
feature is_journal(x:item)
feature is_bell_pepper(x:item)
feature is_shoes(x:item)
feature is_love_seat(x:item)
feature is_facecream(x:item)
feature is_food_bread(x:item)
feature is_cutlery_fork(x:item)
feature is_coffee_pot(x:item)
feature is_pencil(x:item)
feature is_box(x:item)
feature is_sauce(x:item)
feature is_tv(x:item)
feature is_blender(x:item)
feature is_toothbrush(x:item)
feature is_pen(x:item)
feature is_wall(x:item)
feature is_pajamas(x:item)
feature is_spectacles(x:item)
feature is_maindoor(x:item)
feature is_lime(x:item)
feature is_creamybuns(x:item)
feature is_video_game_controller(x:item)
feature is_closetdrawer(x:item)
feature is_instrument_piano(x:item)
feature is_pancake(x:item)
feature is_shirt(x:item)
feature is_laptop(x:item)
feature is_salad(x:item)
feature is_hands_both(x:item)
feature is_conditioner(x:item)
feature is_curtains(x:item)
feature is_pie(x:item)
feature is_candybar(x:item)
feature is_food_vegetable(x:item)
feature is_condiment_bottle(x:item)
feature is_highlighter(x:item)
feature is_pudding(x:item)
feature is_lighting(x:item)
feature is_paper_towel(x:item)
feature is_cupboard(x:item)
feature is_form(x:item)
feature is_clothes_dress(x:item)
feature is_poundcake(x:item)
feature is_food_cake(x:item)
feature is_coffeemaker(x:item)
feature is_board_game(x:item)
feature is_wineglass(x:item)
feature is_kitchen_table(x:item)
feature is_receipt(x:item)
feature is_pants(x:item)
feature is_plum(x:item)
feature is_chips(x:item)
feature is_instrument_guitar(x:item)
feature is_desk(x:item)
feature is_tea_bag(x:item)
feature is_mop_bucket(x:item)
feature is_diary(x:item)
feature is_cupcake(x:item)
feature is_stall(x:item)
feature is_razor(x:item)
feature is_piano_bench(x:item)
feature is_foundation(x:item)
feature is_towel(x:item)
feature is_groceries(x:item)
feature is_legs_both(x:item)
feature is_dining_room(x:item)
feature is_food_cheese(x:item)
feature is_lotionbottle(x:item)
feature is_food_carrots(x:item)
feature is_band_aids(x:item)
feature is_food_onion(x:item)
feature is_floor(x:item)
feature is_dish_bowl(x:item)
feature is_clothes_underwear(x:item)
feature is_mouse_mat(x:item)
feature is_arms_both(x:item)
feature is_woman(x:item)
feature is_rag(x:item)
feature is_toothbrush_holder(x:item)
feature is_soap(x:item)
feature is_ceiling(x:item)
feature is_dry_pasta(x:item)
feature is_computer(x:item)
feature is_bread_slice(x:item)
feature is_cereal(x:item)
feature is_food_fish(x:item)
feature is_crayons(x:item)
feature is_dresser(x:item)
feature is_cup(x:item)
feature is_note_pad(x:item)
feature is_wooden_spoon(x:item)
feature is_food_snack(x:item)
feature is_couch(x:item)
feature is_wall_clock(x:item)
feature is_telephone(x:item)
feature is_lemon(x:item)
feature is_microphone(x:item)
feature is_pantry(x:item)
feature is_food_steak(x:item)
feature is_table(x:item)
feature is_cellphone(x:item)
feature is_electrical_outlet(x:item)
feature is_powersocket(x:item)
feature is_food_banana(x:item)
feature is_teeth(x:item)
feature is_remote_control(x:item)
feature is_hair(x:item)
feature is_alarm_clock(x:item)
feature is_keyboard(x:item)
feature is_food_chicken(x:item)
feature is_doorjamb(x:item)
feature is_home_office(x:item)
feature is_sundae(x:item)
feature is_child(x:item)
feature is_bananas(x:item)
feature is_chessboard(x:item)
feature is_bedroom(x:item)
feature is_dish_soap(x:item)
feature is_crackers(x:item)
feature is_folder(x:item)
feature is_chocolatesyrup(x:item)
feature is_glue(x:item)
feature is_washing_machine(x:item)
feature is_kitchen(x:item)
feature is_after_shave(x:item)
feature is_papertowel(x:item)
feature is_comforter(x:item)
feature is_notebook(x:item)
feature is_placemat(x:item)
feature is_bills(x:item)
feature is_garbage_can(x:item)
feature is_vacuum_cleaner(x:item)
feature is_diningtable(x:item)
feature is_food_apple(x:item)
feature is_door(x:item)
feature is_livingroom(x:item)
feature is_paper(x:item)
feature is_bench(x:item)
feature is_oven(x:item)
feature is_textbook(x:item)
feature is_food_lemon(x:item)
feature is_food_orange(x:item)
feature is_homework(x:item)
feature is_shelf(x:item)
feature is_food_peanut_butter(x:item)



#controllers
controller walk_executor(x: item)
controller switchoff_executor(x: item)
controller switchon_executor(x: item)
controller put_executor(x: item, y: item)
controller putin_executor(x: item, y: item)
controller grab_executor(x: item)
controller standup_executor(x: character)
controller wash_executor(x: item)
controller scrub_executor(x: item)
controller rinse_executor(x: item)
controller sit_executor(x: item)
controller lie_executor(x: item)
controller open_executor(x: item)
controller close_executor(x: item)
controller pour_executor(x: item, y: item)
controller plugin_executor(x: item)
controller plugout_executor(x: item)
controller find_executor(x: item)
controller turnto_executor(x: item)
controller cut_executor(x: item)
controller eat_executor(x: item)
controller sleep_executor(x: character)
controller greet_executor(x: item)
controller drink_executor(x: item)
controller lookat_executor(x: item)
controller wipe_executor(x: item)
controller puton_executor(x: item)
controller putoff_executor(x: item)
controller read_executor(x: item)
controller touch_executor(x: item)
controller type_executor(x: item)
controller watch_executor(x: item)
controller move_executor(x: item)
controller push_executor(x: item)
controller pull_executor(x: item)
controller exp(x:item, y:item)
controller obs(x:item,q:string)
controller echo()

behavior put(inhand_obj: item, obj: item):
  body:
    assert not is_room(obj)
    #assert not pourable(inhand_obj)
    achieve not unknown(obj)
    achieve not unknown(inhand_obj)
    achieve_once inhand(inhand_obj)
    achieve_once close_char(char, obj)
    put_executor(inhand_obj, obj)

  eff:
    holds_rh[char, inhand_obj] = False
    holds_lh[char, inhand_obj] = False
    inhand[inhand_obj] = False
    on[inhand_obj, obj] = True
    close[inhand_obj, obj] = True
    close[obj, inhand_obj] = True
    foreach inter in (findall x: item: close(x, obj) and not unknown(x)):
      close[inter, inhand_obj] = True
      close[inhand_obj, inter] = True
    used[obj] = True
    used[inhand_obj] = True
    has_a_free_hand[char] = True

behavior putin(inhand_obj: item, obj: item):
  body:
    assert recipient(obj) or containers(obj) or can_open(obj) or eatable(obj)
    #assert not pourable(inhand_obj)
    if has_size(obj) and has_size(inhand_obj):
      assert size(inhand_obj) <= size(obj)
    achieve not unknown(obj)
    achieve not unknown(inhand_obj)
    if can_open(obj):
      achieve open(obj)
    achieve_once inhand(inhand_obj)
    achieve_once close_char(char, obj)
    putin_executor(inhand_obj, obj)

  eff:
    holds_rh[char, inhand_obj] = False
    holds_lh[char, inhand_obj] = False
    inhand[inhand_obj] = False
    inside[inhand_obj, obj] = True
    close[inhand_obj, obj] = True
    close[obj, inhand_obj] = True
    foreach inter in (findall x: item: close(x, obj) and not unknown(x)):
      close[inter, inhand_obj] = True
      close[inhand_obj, inter] = True
    foreach inside_obj in (findall x: item: inside(x, inhand_obj)):
      inside[inside_obj, obj] = True
    used[obj] = True
    used[inhand_obj] = True
    has_a_free_hand[char] = True

behavior put_close(inhand_obj: item, obj: item):
  goal: close(inhand_obj, obj)
  body:
    put(inhand_obj, obj)

behavior put_on(inhand_obj: item, obj: item):
  goal: on(inhand_obj, obj)
  body:
    put(inhand_obj, obj)


behavior put_inside(inhand_obj: item, obj: item):
  goal: inside(inhand_obj, obj)
  body:
    putin(inhand_obj, obj)

behavior empty_a_hand(char: character):
  goal: has_a_free_hand(char)
  body:
    assert not has_a_free_hand(char)
    bind surf:item where:
      surfaces(surf)
    bind give_up_obj:item where:
      inhand(give_up_obj)
    put(give_up_obj, surf)
  eff:
    has_a_free_hand[char] = True

behavior stand():
  goal: standing(char)
  body:
    assert sitting(char) or lying(char)
    standup_executor(char)
  eff:
    sitting[char] = False
    lying[char] = False


behavior sit_somewhere(location:item):
  goal: on_char(char, location)
  body:
    assert sittable(location)
    achieve not unknown(location)
    achieve_once close_char(char, location)
    sit_executor(location)
  eff:
    sitting[char] = True
    on_char[char, location] = True
    lying[char] = False

behavior lie_somewhere(location:item):
  goal: on_char(char, location)
  body:
    assert lieable(location)
    achieve not unknown(location)
    achieve_once close_char(char, location)
    lie_executor(location)
  eff:
    lying[char] = True
    sitting[char] = False
    on_char[char, location] = True

def obj_inside_or_on(obj1: item, obj2: item):
  return inside(obj1, obj2) or on(obj2, obj1)

behavior walk_to(obj: item):
  goal: close_char(char, obj)
  body:
    achieve standing(char)
    achieve not unknown(obj)
    walk_executor(obj)
    let inhand_objects=findall o: item where: inhand(o)

  eff:
    inside_char[char, :] = False
    close_char[char, :] = False
    facing_char[char, :] = False
    foreach o in inhand_objects:
      inside[o, :]= False
      close[o, :] = False
      close[:, o] = False

    foreach icf in (findall t:item: obj_inside_or_on(obj, t)):
      close_char[char, icf] = True
      if not (can_open(icf) and closed(icf)):
        unknown[icf] = False
      foreach o in inhand_objects:
        close[o, icf] = True
        close[icf, o] = True

    close_char[char,obj] = True
    foreach o in inhand_objects:
      close[o, obj] = True
      close[obj, o] = True

behavior find(obj:item):
  goal: facing_char(char, obj) and close_char(char, obj)
  body:
    achieve not unknown(obj)
    if on_body(obj, char):
      find_executor(obj)
    else:
      achieve_once close_char(char, obj)
      find_executor(obj)
  eff:
    foreach o in (findall t:item: facing_char(char, t)):
      facing_char[char, o] = False
    facing_char[char, obj] = True

behavior turnto(obj:item):
  goal: facing_char(char, obj)
  body:
    achieve not unknown(obj)
    turnto_executor(obj)
  eff:
    foreach o in (findall t:item: facing_char(char, t)):
      facing_char[char, o] = False
    facing_char[char, obj] = True

behavior switch_off(obj: item):
  goal: is_off(obj)
  body:
    assert has_switch(obj)
    achieve not unknown(obj)
    achieve_once has_a_free_hand(char)
    achieve_once close_char(char, obj)
    switchoff_executor(obj)
  eff:
    is_off[obj] = True
    is_on[obj] = False
    used[obj] = True

behavior switch_on(obj: item):
  goal: is_on(obj)
  body:
    assert has_switch(obj)
    achieve_once has_a_free_hand(char)
    achieve not unknown(obj)
    if has_plug(obj):
      achieve plugged(obj)
    if can_open(obj) and not is_stove(obj):
      achieve closed(obj)
    achieve_once close_char(char, obj)
    switchon_executor(obj)
  eff:
    is_off[obj] = False
    is_on[obj] = True
    used[obj] = True

behavior grab(obj: item):
  goal: inhand(obj)
  body:
    assert grabbable(obj) or is_water(obj)
    achieve not unknown(obj)
    achieve_once has_a_free_hand(char)
    foreach obj2:item:
      if inside(obj,obj2) and can_open(obj2):
          achieve_once open(obj2)
    achieve_once close_char(char, obj)
    grab_executor(obj)
  eff:
    inhand[obj] = True
    on[obj, :] = False
    inside[obj, :] = False
    close[obj, :] = False
    close[:, obj] = False
    if exists item1: item : holds_lh(char, item1):
      holds_rh[char, obj] = True
      has_a_free_hand[char] = False
    else:
      holds_lh[char, obj] = True
    close_char[char,obj]=True
    used[obj] = True

#behavior wash(obj: item):
#  goal: clean(obj)
#  body:
#    assert grabbable(obj) or is_water(obj)
#    achieve not unknown(obj)
#    achieve_once has_a_free_hand(char)
#    achieve_once close_char(char, obj)
#    wash_executor(obj)
#  eff:
#    dirty[obj] = False
#    clean[obj] = True
#    used[obj] = True

behavior wash(obj: item):
  goal: clean(obj)
  body:
    achieve not unknown(obj)
    symbol obj_inside_sink=exists sink:item: is_sink(sink) and inside(obj, sink)
    if not obj_inside_sink:
      bind sink:item where:
        is_sink(sink)
      achieve_once inside(obj, sink)
    wash_executor(obj)
  eff:
    dirty[obj] = False
    clean[obj] = True
    used[obj] = True

behavior scrub(obj: item):
  body:
    achieve not unknown(obj)
    achieve_once has_a_free_hand(char)
    achieve_once close_char(char, obj)
    scrub_executor(obj)
  eff:
    dirty[obj] = False
    clean[obj] = True
    used[obj] = True

behavior rinse(obj: item):
  body:
    achieve not unknown(obj)
    achieve_once has_a_free_hand(char)
    achieve_once close_char(char, obj)
    rinse_executor(obj)
  eff:
    dirty[obj] = False
    clean[obj] = True
    used[obj] = True

behavior opens(obj: item):
  goal: open(obj)
  body:
    assert can_open(obj)
    achieve not unknown(obj)
    achieve_once has_a_free_hand(char)
    if has_switch(obj) and is_on(obj):
      achieve is_off(obj)
    achieve_once close_char(char, obj)
    symbol containers=exists item1:item: inside(obj, item1) and can_open(item1)
    if containers:
      bind container:item where:
        inside(obj, container) and can_open(container)
      achieve open(container)
    open_executor(obj)
  eff:
    open[obj] = True
    closed[obj] = False
    foreach i in (findall x: item: inside(x, obj)):
      unknown[i] = False
    used[obj] = True

behavior closes(obj: item):
  goal: closed(obj)
  body:
    assert can_open(obj)
    achieve not unknown(obj)
    achieve_once has_a_free_hand(char)
    achieve_once close_char(char, obj)
    close_executor(obj)
  eff:
    open[obj] = False
    closed[obj] = True
    used[obj] = True

#def pour_target(obj: item):
#  return is_hands_both(obj) or is_sponge(obj) or is_face(obj)

#behavior pour_in(obj: item, target: item):
#  goal: inside(obj, target)
#  body:
#    assert (pourable(obj) or drinkable(obj)) and recipient(target)
#    assert recipient(target) or pour_target(obj)
#    achieve not unknown(obj)
#    achieve not unknown(target)
#    achieve inhand(obj)
#    achieve close_char(char, target)
#    pour_executor(obj, target)
#  eff:
#    inside[obj, target] = True
#    if is_water(obj):
#      holds_lh[char, obj] = False
#      holds_rh[char, obj] = False

#behavior pour_on(obj: item, target: item):
#  goal: inside(obj, target)
#  body:
#    assert (pourable(obj) or drinkable(obj)) and recipient(target)
#    achieve not unknown(obj)
#    achieve not unknown(target)
#    achieve inhand(obj)
#    achieve close_char(char, target)
#    pour_executor(obj, target)
#  eff:
#    on[obj, target] = True
#    if is_water(obj):
#      holds_lh[char, obj] = False
#      holds_rh[char, obj] = False

behavior plugin(object:item):
  goal: plugged(object)
  body:
    assert has_plug(object)
    achieve not unknown(object)
    achieve_once has_a_free_hand(char)
    achieve_once close_char(char, object)
    plugin_executor(object)
  eff:
    plugged[object] = True
    unplugged[object] = False
    used[object] = True

behavior plugout(object:item):
  goal: unplugged(object)
  body:
    assert has_plug(object)
    achieve not unknown(object)
    achieve_once has_a_free_hand(char)
    if has_switch(object):
      achieve is_off(object)
    achieve_once close_char(char, object)
    plugout_executor(object)
  eff:
    plugged[object] = False
    unplugged[object] = True
    used[object] = True

behavior cuts(object:item):
  goal: cut(object)
  body:
    assert cuttable(object) or eatable(object)
    achieve not unknown(object)
    symbol has_cutting_board=exists item1:item: is_cutting_board(item1)
    if has_cutting_board:
      bind cutting_board:item where:
        is_cutting_board(cutting_board)
      achieve_once on(object, cutting_board)
    symbol has_knife=exists knife:item: is_knife(knife) and inhand(knife)
    if not has_knife:
      bind new_knife:item where:
        is_knife(new_knife)
      achieve_once inhand(new_knife)
    achieve_once close_char(char, object)
    cut_executor(object)
  eff:
    cut[object] = True
    used[object] = True

behavior eat(object:item):
  body:
    assert eatable(object)
    achieve not unknown(object)
    eat_executor(object)
  eff:
    used[object] = True


behavior sleep_somewhere(location:item):
  body:
    symbol has_lieable_place=exists item1:item: lieable(item1)
    symbol has_sittable_place=exists item2:item: sittable(item2)
    assert has_lieable_place or has_sittable_place
    if has_lieable_place:
      lie_somewhere(location)
    else:
      sit_somewhere(location)
  eff:
    sleeping[char] = True

behavior wake_up():
  goal: not sleeping(char)
  body:
    assert sleeping(char)
    stand()
  eff:
    sleeping[char] = False

behavior wipe(obj:item):
  body:
    symbol has_cleaning_solution=exists item1:item: is_towel(item1) or is_rag(item1) or is_sponge(item1) or is_paper_towel(item1) or is_cloth_napkin(item1) or is_duster(item1) or is_cleaning_solution(item1)
    if not has_cleaning_solution:
      bind cleaning_tool:item where:
        is_towel(cleaning_tool) or is_rag(cleaning_tool) or is_sponge(cleaning_tool) or is_paper_towel(cleaning_tool) or is_cloth_napkin(cleaning_tool) or is_duster(cleaning_tool) or is_cleaning_solution(cleaning_tool)
      achieve not unknown(cleaning_tool)
      achieve_once inhand(cleaning_tool)
    achieve_once close_char(char, obj)
    wipe_executor(obj)
  eff:
    dirty[obj] = False
    clean[obj] = True
    used[obj] = True

behavior put_on_body(inhand_obj: item):
  goal: on_body(inhand_obj, char)
  body:
    assert is_clothes(inhand_obj)
    achieve not unknown(inhand_obj)
    achieve_once inhand(inhand_obj)
    puton_executor(inhand_obj)
  eff:
    on_body[inhand_obj, char] = True
    used[inhand_obj] = True

behavior put_off_body(clo: item):
  goal: not on_body(clo, char)
  body:
    assert is_clothes(clo)
    putoff_executor(clo)
  eff:
    on_body[clo, char] = False
    used[clo] = True

behavior get_water(obj:item):
  goal: has_water(obj)
  body:
    symbol has_faucet_around=exists faucet:item: is_faucet(faucet) and close(obj, faucet)
    if grabbable(obj):
      bind faucet:item where:
        is_faucet(faucet)
      if can_open(obj):
        achieve open(obj)
      achieve inhand(obj)
      achieve_once close_char(char, faucet)
      achieve_once is_on(faucet)
      achieve_once is_off(faucet)
    else:
      if has_faucet_around:
        bind faucet:item where:
          is_faucet(faucet) and close(obj, faucet)
        achieve_once is_on(faucet)
        achieve_once is_off(faucet)
  eff:
    has_water[obj] = True

behavior read(material:item):
  body:
    assert readable(material)
    achieve not unknown(material)
    achieve inhand(material)
    read_executor(material)
  eff:
    used[material] = True

behavior touch(obj:item):
  body:
    achieve not unknown(obj)
    foreach obj2:item:
      if inside(obj,obj2):
        if not is_room(obj2):
          assert can_open(obj2) or recipient(obj2) or eatable(obj2)
          if can_open(obj2):
            achieve open(obj2)
    achieve_once close_char(char, obj)
    touch_executor(obj)
  eff:
    used[obj] = True

behavior type(obj:item):
  body:
    assert is_keyboard(obj) or has_switch(obj)
    achieve not unknown(obj)

    achieve close_char(char, obj)
    type_executor(obj)
  eff:
    used[obj] = True

behavior watch(obj:item):
  body:
    assert lookable(obj)
    achieve not unknown(obj)
    achieve facing_char(char, obj)
  eff:
    used[obj] = True

behavior drink(obj: item):
  body:
    assert drinkable(obj) or recipient(obj)
    achieve not unknown(obj)
    achieve_once inhand(obj)
    drink_executor(obj)
  eff:
    used[obj] = True

behavior look_at(obj:item):
  body:
    achieve not unknown(obj)
    achieve_once facing_char(char, obj)
    lookat_executor(obj)
  eff:
    used[obj] = True

behavior greet(person:item):
  body:
    assert person(person)
    achieve not unknown(person)
    greet_executor(person)
  eff:
    used[person] = True

behavior move(obj:item):
  body:
    assert movable(obj) or is_button(obj) or is_chair(obj) or is_curtain(obj)
    achieve not unknown(obj)
    achieve_once has_a_free_hand(char)
    achieve_once close_char(char, obj)
    move_executor(obj)
  eff:
    used[obj] = True

behavior push(obj:item):
  body:
    assert movable(obj) or is_button(obj) or is_chair(obj) or is_curtain(obj)
    achieve not unknown(obj)
    achieve_once has_a_free_hand(char)
    achieve_once close_char(char, obj)
    push_executor(obj)
  eff:
    used[obj] = True

behavior pull(obj:item):
  body:
    assert movable(obj) or is_button(obj) or is_chair(obj) or is_curtain(obj)
    achieve not unknown(obj)
    achieve_once has_a_free_hand(char)
    achieve_once close_char(char, obj)
    pull_executor(obj)
  eff:
    used[obj] = True

behavior squeeze(obj:item):
  body:
    assert is_cleaning_solution(obj) or is_tooth_paste(obj) or is_shampoo(obj) or is_dish_soap(obj) or is_soap(obj) or is_towel(obj) or is_rag(obj) or has_paper(obj) or is_sponge(obj) or is_food_lemon(obj) or is_clothes(obj) or is_check(obj)
    achieve not unknown(obj)
    achieve_once has_a_free_hand(char)
    achieve_once close_char(char, obj)
  eff:
    used[obj] = True

behavior observe(obj:item, q:string):
  body:
    achieve not unknown(obj)
    achieve_once close_char(char, obj)
    if can_open(obj):
      achieve_once open(obj)
    obs(obj,q)
  eff:
    visited[obj] = True

behavior visit(item:item):
  goal: visited(item)
  body:
    observe(item,"look around this place")
