problem "agent-problem"
domain "virtualhome_partial.cdl"

#!pragma planner_is_goal_serializable=False
#!pragma planner_is_goal_ordered=True
#!pragma planner_always_commit_skeleton=True

objects:
#objects
  clothes_pants_2085:item
  clothes_shirt_2086:item
  clothes_socks_2087:item
  clothes_skirt_2088:item
  iron_2089:item
  basket_for_clothes_2006:item
  washing_machine_2007:item
  food_steak_2008:item
  food_apple_2009:item
  food_bacon_2010:item
  food_banana_2011:item
  food_bread_2012:item
  food_cake_2013:item
  food_carrot_2014:item
  food_cereal_2015:item
  food_cheese_2016:item
  food_chicken_2017:item
  food_dessert_2018:item
  food_donut_2019:item
  food_egg_2020:item
  food_fish_2021:item
  food_food_2022:item
  food_fruit_2023:item
  food_hamburger_2024:item
  food_ice_cream_2025:item
  food_jam_2026:item
  food_kiwi_2027:item
  food_lemon_2028:item
  food_noodles_2029:item
  food_oatmeal_2030:item
  food_orange_2031:item
  food_onion_2032:item
  food_peanut_butter_2033:item
  food_pizza_2034:item
  food_potato_2035:item
  food_rice_2036:item
  food_salt_2037:item
  food_snack_2038:item
  food_sugar_2039:item
  food_turkey_2040:item
  food_vegetable_2041:item
  dry_pasta_2042:item
  milk_2043:item
  clothes_dress_2044:item
  clothes_hat_2045:item
  clothes_gloves_2046:item
  clothes_jacket_2047:item
  clothes_scarf_2048:item
  clothes_underwear_2049:item
  knife_2050:item
  cutting_board_2051:item
  remote_control_2052:item
  soap_2053:item
  soap_2054:item
  cat_2055:item
  towel_2056:item
  towel_2057:item
  towel_2058:item
  towel_2059:item
  cd_player_2060:item
  dvd_player_2061:item
  headset_2062:item
  cup_2063:item
  cup_2064:item
  stove_2065:item
  book_2066:item
  book_2067:item
  coffee_table_2068:item
  pot_2069:item
  vacuum_cleaner_2070:item
  bowl_2071:item
  bowl_2072:item
  cleaning_solution_2073:item
  ironing_board_2074:item
  cd_2075:item
  headset_2076:item
  phone_2077:item
  sauce_2078:item
  oil_2079:item
  fork_2080:item
  fork_2081:item
  spectacles_2082:item
  fryingpan_2083:item
  detergent_2084:item
  bathroom_1:item
  floor_2:item
  floor_3:item
  floor_4:item
  floor_5:item
  floor_6:item
  floor_7:item
  floor_8:item
  wall_9:item
  wall_10:item
  wall_11:item
  wall_12:item
  wall_13:item
  wall_14:item
  wall_15:item
  ceiling_16:item
  ceiling_17:item
  ceiling_18:item
  ceiling_19:item
  ceiling_20:item
  ceiling_21:item
  mat_22:item
  curtain_23:item
  curtain_24:item
  curtain_25:item
  ceilinglamp_26:item
  walllamp_27:item
  walllamp_28:item
  walllamp_29:item
  bathtub_30:item
  towel_rack_31:item
  towel_rack_32:item
  towel_rack_33:item
  towel_rack_34:item
  wallshelf_35:item
  shower_36:item
  toilet_37:item
  shower_38:item
  curtain_39:item
  bathroom_cabinet_40:item
  bathroom_counter_41:item
  sink_42:item
  faucet_43:item
  door_44:item
  doorjamb_45:item
  window_63:item
  light_64:item
  bedroom_67:item
  floor_68:item
  floor_69:item
  floor_70:item
  floor_71:item
  floor_72:item
  floor_73:item
  floor_74:item
  floor_75:item
  floor_76:item
  floor_77:item
  wall_78:item
  wall_79:item
  wall_80:item
  wall_81:item
  wall_82:item
  wall_83:item
  wall_84:item
  wall_85:item
  window_86:item
  ceiling_87:item
  ceiling_88:item
  ceiling_89:item
  ceiling_90:item
  ceiling_91:item
  ceiling_92:item
  ceiling_93:item
  ceiling_94:item
  ceiling_95:item
  ceilinglamp_96:item
  tablelamp_97:item
  tablelamp_98:item
  trashcan_99:item
  nightstand_100:item
  bookshelf_101:item
  nightstand_102:item
  chair_103:item
  desk_104:item
  bed_105:item
  chair_106:item
  table_107:item
  dresser_108:item
  hanger_109:item
  hanger_110:item
  hanger_111:item
  hanger_112:item
  hanger_113:item
  hanger_114:item
  hanger_115:item
  closetdrawer_116:item
  closetdrawer_117:item
  closetdrawer_118:item
  closetdrawer_119:item
  closetdrawer_120:item
  closetdrawer_121:item
  closetdrawer_122:item
  dresser_123:item
  hanger_124:item
  hanger_126:item
  hanger_128:item
  hanger_130:item
  hanger_132:item
  hanger_134:item
  hanger_136:item
  hanger_138:item
  hanger_140:item
  hanger_141:item
  hanger_142:item
  closetdrawer_143:item
  closetdrawer_146:item
  closetdrawer_148:item
  closetdrawer_150:item
  closetdrawer_154:item
  closetdrawer_158:item
  closetdrawer_160:item
  doorjamb_165:item
  mouse_166:item
  mousepad_167:item
  keyboard_168:item
  light_169:item
  computer_170:item
  cpuscreen_171:item
  mat_173:item
  drawing_174:item
  drawing_175:item
  drawing_176:item
  orchid_178:item
  curtain_179:item
  curtain_180:item
  curtain_181:item
  pillow_182:item
  pillow_183:item
  photoframe_185:item
  dining_room_201:item
  floor_202:item
  floor_203:item
  floor_204:item
  floor_205:item
  floor_206:item
  floor_207:item
  floor_208:item
  wall_209:item
  wall_210:item
  wall_211:item
  wall_212:item
  wall_213:item
  wall_214:item
  wall_215:item
  ceiling_216:item
  ceiling_217:item
  ceiling_218:item
  ceiling_219:item
  ceiling_220:item
  ceiling_221:item
  door_222:item
  ceilinglamp_223:item
  ceilinglamp_224:item
  tvstand_225:item
  table_226:item
  bench_227:item
  bench_228:item
  cupboard_229:item
  kitchen_counter_230:item
  sink_231:item
  faucet_232:item
  bookshelf_233:item
  wallshelf_234:item
  wallshelf_235:item
  mat_236:item
  mat_237:item
  drawing_238:item
  drawing_239:item
  drawing_240:item
  drawing_241:item
  drawing_242:item
  drawing_243:item
  orchid_244:item
  light_245:item
  powersocket_246:item
  phone_247:item
  television_248:item
  wall_clock_249:item
  photoframe_285:item
  stovefan_288:item
  fridge_289:item
  coffe_maker_290:item
  toaster_292:item
  oven_295:item
  tray_296:item
  microwave_297:item
  home_office_319:item
  floor_320:item
  floor_321:item
  floor_322:item
  floor_323:item
  floor_324:item
  floor_325:item
  floor_326:item
  floor_327:item
  floor_328:item
  wall_329:item
  wall_330:item
  wall_331:item
  wall_332:item
  wall_333:item
  wall_334:item
  wall_335:item
  wall_336:item
  ceiling_337:item
  ceiling_338:item
  ceiling_339:item
  ceiling_340:item
  ceiling_341:item
  ceiling_342:item
  ceiling_343:item
  ceiling_344:item
  ceiling_345:item
  doorjamb_346:item
  doorjamb_347:item
  window_348:item
  ceilinglamp_349:item
  walllamp_350:item
  walllamp_351:item
  couch_352:item
  tvstand_353:item
  bookshelf_354:item
  table_355:item
  chair_356:item
  desk_357:item
  dresser_358:item
  hanger_359:item
  hanger_361:item
  hanger_363:item
  hanger_365:item
  hanger_367:item
  hanger_369:item
  hanger_372:item
  hanger_374:item
  hanger_375:item
  hanger_376:item
  closetdrawer_377:item
  closetdrawer_380:item
  closetdrawer_382:item
  closetdrawer_384:item
  closetdrawer_388:item
  closetdrawer_392:item
  closetdrawer_394:item
  filing_cabinet_399:item
  drawing_400:item
  mat_401:item
  drawing_402:item
  drawing_403:item
  drawing_404:item
  pillow_405:item
  pillow_406:item
  curtain_407:item
  curtain_408:item
  curtain_409:item
  television_410:item
  light_411:item
  powersocket_412:item
  mouse_413:item
  mousepad_414:item
  keyboard_415:item
  cpuscreen_416:item
  computer_417:item
  photoframe_430:item
  plate_1000:item
  dishwasher_1001:item
  coffee_filter_2000:item
  pencil_2001:item
  hairbrush_2002:item
  drawing_2003:item
  chair_2004:item
  napkin_2005:item
#object_end

init:
    #categories
    is_pants[clothes_pants_2085]=True
    is_clothes_pants[clothes_pants_2085]=True
    is_shirt[clothes_shirt_2086]=True
    is_clothes_shirt[clothes_shirt_2086]=True
    is_clothes_socks[clothes_socks_2087]=True
    is_clothes_skirt[clothes_skirt_2088]=True
    is_iron[iron_2089]=True
    is_clothes_pile[basket_for_clothes_2006]=True
    is_basket_for_clothes[basket_for_clothes_2006]=True
    is_washing_machine[washing_machine_2007]=True
    is_food_steak[food_steak_2008]=True
    is_food_apple[food_apple_2009]=True
    is_apple[food_apple_2009]=True
    is_food_bacon[food_bacon_2010]=True
    is_banana[food_banana_2011]=True
    is_food_banana[food_banana_2011]=True
    is_bread_slice[food_bread_2012]=True
    is_bread[food_bread_2012]=True
    is_food_bread[food_bread_2012]=True
    is_food_cake[food_cake_2013]=True
    is_carrot[food_carrot_2014]=True
    is_food_carrot[food_carrot_2014]=True
    is_food_cereal[food_cereal_2015]=True
    is_cereal[food_cereal_2015]=True
    is_food_cheese[food_cheese_2016]=True
    is_food_chicken[food_chicken_2017]=True
    is_chicken[food_chicken_2017]=True
    is_watermelon[food_dessert_2018]=True
    is_poundcake[food_dessert_2018]=True
    is_milkshake[food_dessert_2018]=True
    is_sundae[food_dessert_2018]=True
    is_food_dessert[food_dessert_2018]=True
    is_creamybuns[food_dessert_2018]=True
    is_pudding[food_dessert_2018]=True
    is_pie[food_dessert_2018]=True
    is_pancake[food_dessert_2018]=True
    is_cupcake[food_dessert_2018]=True
    is_food_donut[food_donut_2019]=True
    is_food_egg[food_egg_2020]=True
    is_food_fish[food_fish_2021]=True
    is_salmon[food_fish_2021]=True
    is_pear[food_food_2022]=True
    is_salmon[food_food_2022]=True
    is_creamybuns[food_food_2022]=True
    is_whippedcream[food_food_2022]=True
    is_orange[food_food_2022]=True
    is_food_food[food_food_2022]=True
    is_bell_pepper[food_food_2022]=True
    is_cutlets[food_food_2022]=True
    is_cucumber[food_food_2022]=True
    is_tomato[food_food_2022]=True
    is_bananas[food_food_2022]=True
    is_crackers[food_food_2022]=True
    is_cereal[food_food_2022]=True
    is_chicken[food_food_2022]=True
    is_apple[food_food_2022]=True
    is_bellpepper[food_food_2022]=True
    is_plum[food_food_2022]=True
    is_banana[food_food_2022]=True
    is_chocolatesyrup[food_food_2022]=True
    is_chinesefood[food_food_2022]=True
    is_potato[food_food_2022]=True
    is_pear[food_fruit_2023]=True
    is_plum[food_fruit_2023]=True
    is_watermelon[food_fruit_2023]=True
    is_banana[food_fruit_2023]=True
    is_food_fruit[food_fruit_2023]=True
    is_apple[food_fruit_2023]=True
    is_orange[food_fruit_2023]=True
    is_food_hamburger[food_hamburger_2024]=True
    is_mincedmeat[food_hamburger_2024]=True
    is_food_ice_cream[food_ice_cream_2025]=True
    is_food_jam[food_jam_2026]=True
    is_food_kiwi[food_kiwi_2027]=True
    is_food_lemon[food_lemon_2028]=True
    is_lemon[food_lemon_2028]=True
    is_food_noodles[food_noodles_2029]=True
    is_food_oatmeal[food_oatmeal_2030]=True
    is_cereal[food_oatmeal_2030]=True
    is_food_orange[food_orange_2031]=True
    is_food_onion[food_onion_2032]=True
    is_food_peanut_butter[food_peanut_butter_2033]=True
    is_food_pizza[food_pizza_2034]=True
    is_potato[food_potato_2035]=True
    is_food_potato[food_potato_2035]=True
    is_food_rice[food_rice_2036]=True
    is_condiment_shaker[food_salt_2037]=True
    is_food_salt[food_salt_2037]=True
    is_crackers[food_snack_2038]=True
    is_salt_crackers[food_snack_2038]=True
    is_chips[food_snack_2038]=True
    is_banana[food_snack_2038]=True
    is_candybar[food_snack_2038]=True
    is_apple[food_snack_2038]=True
    is_cupcake[food_snack_2038]=True
    is_food_snack[food_snack_2038]=True
    is_poundcake[food_snack_2038]=True
    is_condiment_shaker[food_sugar_2039]=True
    is_food_sugar[food_sugar_2039]=True
    is_chicken[food_turkey_2040]=True
    is_food_turkey[food_turkey_2040]=True
    is_food_vegetable[food_vegetable_2041]=True
    is_cucumber[food_vegetable_2041]=True
    is_tomato[food_vegetable_2041]=True
    is_carrot[food_vegetable_2041]=True
    is_potato[food_vegetable_2041]=True
    is_salad[food_vegetable_2041]=True
    is_dry_pasta[dry_pasta_2042]=True
    is_milk[milk_2043]=True
    is_clothes_dress[clothes_dress_2044]=True
    is_clothes_hat[clothes_hat_2045]=True
    is_clothes_gloves[clothes_gloves_2046]=True
    is_clothes_jacket[clothes_jacket_2047]=True
    is_clothes_scarf[clothes_scarf_2048]=True
    is_clothes_underwear[clothes_underwear_2049]=True
    is_cutlery_knife[knife_2050]=True
    is_knife[knife_2050]=True
    is_chefknife[knife_2050]=True
    is_cutting_board[cutting_board_2051]=True
    is_controller[remote_control_2052]=True
    is_remote_control[remote_control_2052]=True
    is_soap[soap_2053]=True
    is_barsoap[soap_2053]=True
    is_soap[soap_2054]=True
    is_barsoap[soap_2054]=True
    is_cat[cat_2055]=True
    is_towel[towel_2056]=True
    is_towel[towel_2057]=True
    is_towel[towel_2058]=True
    is_towel[towel_2059]=True
    is_cd_player[cd_player_2060]=True
    is_radio[cd_player_2060]=True
    is_dvd_player[dvd_player_2061]=True
    is_headset[headset_2062]=True
    is_mug[cup_2063]=True
    is_waterglass[cup_2063]=True
    is_wineglass[cup_2063]=True
    is_cup[cup_2063]=True
    is_mug[cup_2064]=True
    is_waterglass[cup_2064]=True
    is_wineglass[cup_2064]=True
    is_cup[cup_2064]=True
    is_stove[stove_2065]=True
    is_oven[stove_2065]=True
    is_textbook[book_2066]=True
    is_novel[book_2066]=True
    is_book[book_2066]=True
    is_textbook[book_2067]=True
    is_novel[book_2067]=True
    is_book[book_2067]=True
    is_kitchen_table[coffee_table_2068]=True
    is_coffeetable[coffee_table_2068]=True
    is_table[coffee_table_2068]=True
    is_diningtable[coffee_table_2068]=True
    is_coffee_table[coffee_table_2068]=True
    is_pot[pot_2069]=True
    is_vacuum_cleaner[vacuum_cleaner_2070]=True
    is_dish_bowl[bowl_2071]=True
    is_bowl[bowl_2071]=True
    is_dish_bowl[bowl_2072]=True
    is_bowl[bowl_2072]=True
    is_cleaning_solution[cleaning_solution_2073]=True
    is_dishwashingliquid[cleaning_solution_2073]=True
    is_ironing_board[ironing_board_2074]=True
    is_cd[cd_2075]=True
    is_headset[headset_2076]=True
    is_wall_phone[phone_2077]=True
    is_phone[phone_2077]=True
    is_cellphone[phone_2077]=True
    is_condiment_bottle[sauce_2078]=True
    is_sauce[sauce_2078]=True
    is_oil[oil_2079]=True
    is_condiment_bottle[oil_2079]=True
    is_fork[fork_2080]=True
    is_cutlery_fork[fork_2080]=True
    is_fork[fork_2081]=True
    is_cutlery_fork[fork_2081]=True
    is_glasses[spectacles_2082]=True
    is_spectacles[spectacles_2082]=True
    is_fryingpan[fryingpan_2083]=True
    is_detergent[detergent_2084]=True
    is_dishwashingliquid[detergent_2084]=True
    is_bathroom[bathroom_1]=True
    is_floor[floor_2]=True
    is_floor[floor_3]=True
    is_floor[floor_4]=True
    is_floor[floor_5]=True
    is_floor[floor_6]=True
    is_floor[floor_7]=True
    is_floor[floor_8]=True
    is_wall[wall_9]=True
    is_wall[wall_10]=True
    is_wall[wall_11]=True
    is_wall[wall_12]=True
    is_wall[wall_13]=True
    is_wall[wall_14]=True
    is_wall[wall_15]=True
    is_ceiling[ceiling_16]=True
    is_ceiling[ceiling_17]=True
    is_ceiling[ceiling_18]=True
    is_ceiling[ceiling_19]=True
    is_ceiling[ceiling_20]=True
    is_ceiling[ceiling_21]=True
    is_rug[mat_22]=True
    is_mat[mat_22]=True
    is_curtain[curtain_23]=True
    is_curtains[curtain_23]=True
    is_curtain[curtain_24]=True
    is_curtains[curtain_24]=True
    is_curtain[curtain_25]=True
    is_curtains[curtain_25]=True
    is_ceilinglamp[ceilinglamp_26]=True
    is_walllamp[walllamp_27]=True
    is_walllamp[walllamp_28]=True
    is_walllamp[walllamp_29]=True
    is_bathtub[bathtub_30]=True
    is_towel_rack[towel_rack_31]=True
    is_towel_rack[towel_rack_32]=True
    is_towel_rack[towel_rack_33]=True
    is_towel_rack[towel_rack_34]=True
    is_wallshelf[wallshelf_35]=True
    is_stall[shower_36]=True
    is_shower[shower_36]=True
    is_toilet[toilet_37]=True
    is_stall[shower_38]=True
    is_shower[shower_38]=True
    is_curtain[curtain_39]=True
    is_curtains[curtain_39]=True
    is_bathroom_cabinet[bathroom_cabinet_40]=True
    is_bathroom_counter[bathroom_counter_41]=True
    is_sink[sink_42]=True
    is_faucet[faucet_43]=True
    is_door[door_44]=True
    is_doorjamb[doorjamb_45]=True
    is_window[window_63]=True
    is_light_switch[light_64]=True
    is_lightswitch[light_64]=True
    is_light[light_64]=True
    is_bedroom[bedroom_67]=True
    is_floor[floor_68]=True
    is_floor[floor_69]=True
    is_floor[floor_70]=True
    is_floor[floor_71]=True
    is_floor[floor_72]=True
    is_floor[floor_73]=True
    is_floor[floor_74]=True
    is_floor[floor_75]=True
    is_floor[floor_76]=True
    is_floor[floor_77]=True
    is_wall[wall_78]=True
    is_wall[wall_79]=True
    is_wall[wall_80]=True
    is_wall[wall_81]=True
    is_wall[wall_82]=True
    is_wall[wall_83]=True
    is_wall[wall_84]=True
    is_wall[wall_85]=True
    is_window[window_86]=True
    is_ceiling[ceiling_87]=True
    is_ceiling[ceiling_88]=True
    is_ceiling[ceiling_89]=True
    is_ceiling[ceiling_90]=True
    is_ceiling[ceiling_91]=True
    is_ceiling[ceiling_92]=True
    is_ceiling[ceiling_93]=True
    is_ceiling[ceiling_94]=True
    is_ceiling[ceiling_95]=True
    is_ceilinglamp[ceilinglamp_96]=True
    is_tablelamp[tablelamp_97]=True
    is_tablelamp[tablelamp_98]=True
    is_garbage_can[trashcan_99]=True
    is_trashcan[trashcan_99]=True
    is_nightstand[nightstand_100]=True
    is_bookshelf[bookshelf_101]=True
    is_nightstand[nightstand_102]=True
    is_chair[chair_103]=True
    is_desk[desk_104]=True
    is_cpu_table[desk_104]=True
    is_bed[bed_105]=True
    is_chair[chair_106]=True
    is_coffee_table[table_107]=True
    is_kitchen_table[table_107]=True
    is_table[table_107]=True
    is_diningtable[table_107]=True
    is_closet[dresser_108]=True
    is_dresser[dresser_108]=True
    is_coatrack[hanger_109]=True
    is_hanger[hanger_109]=True
    is_coatrack[hanger_110]=True
    is_hanger[hanger_110]=True
    is_coatrack[hanger_111]=True
    is_hanger[hanger_111]=True
    is_coatrack[hanger_112]=True
    is_hanger[hanger_112]=True
    is_coatrack[hanger_113]=True
    is_hanger[hanger_113]=True
    is_coatrack[hanger_114]=True
    is_hanger[hanger_114]=True
    is_coatrack[hanger_115]=True
    is_hanger[hanger_115]=True
    is_closetdrawer[closetdrawer_116]=True
    is_closetdrawer[closetdrawer_117]=True
    is_closetdrawer[closetdrawer_118]=True
    is_closetdrawer[closetdrawer_119]=True
    is_closetdrawer[closetdrawer_120]=True
    is_closetdrawer[closetdrawer_121]=True
    is_closetdrawer[closetdrawer_122]=True
    is_closet[dresser_123]=True
    is_dresser[dresser_123]=True
    is_coatrack[hanger_124]=True
    is_hanger[hanger_124]=True
    is_coatrack[hanger_126]=True
    is_hanger[hanger_126]=True
    is_coatrack[hanger_128]=True
    is_hanger[hanger_128]=True
    is_coatrack[hanger_130]=True
    is_hanger[hanger_130]=True
    is_coatrack[hanger_132]=True
    is_hanger[hanger_132]=True
    is_coatrack[hanger_134]=True
    is_hanger[hanger_134]=True
    is_coatrack[hanger_136]=True
    is_hanger[hanger_136]=True
    is_coatrack[hanger_138]=True
    is_hanger[hanger_138]=True
    is_coatrack[hanger_140]=True
    is_hanger[hanger_140]=True
    is_coatrack[hanger_141]=True
    is_hanger[hanger_141]=True
    is_coatrack[hanger_142]=True
    is_hanger[hanger_142]=True
    is_closetdrawer[closetdrawer_143]=True
    is_closetdrawer[closetdrawer_146]=True
    is_closetdrawer[closetdrawer_148]=True
    is_closetdrawer[closetdrawer_150]=True
    is_closetdrawer[closetdrawer_154]=True
    is_closetdrawer[closetdrawer_158]=True
    is_closetdrawer[closetdrawer_160]=True
    is_doorjamb[doorjamb_165]=True
    is_mouse[mouse_166]=True
    is_mouse_mat[mousepad_167]=True
    is_mousemat[mousepad_167]=True
    is_mousepad[mousepad_167]=True
    is_keyboard[keyboard_168]=True
    is_light_switch[light_169]=True
    is_lightswitch[light_169]=True
    is_light[light_169]=True
    is_cpu_case[computer_170]=True
    is_pc[computer_170]=True
    is_computer[computer_170]=True
    is_cpuscreen[cpuscreen_171]=True
    is_rug[mat_173]=True
    is_mat[mat_173]=True
    is_wallpictureframe[drawing_174]=True
    is_drawing[drawing_174]=True
    is_wallpictureframe[drawing_175]=True
    is_drawing[drawing_175]=True
    is_wallpictureframe[drawing_176]=True
    is_drawing[drawing_176]=True
    is_orchid[orchid_178]=True
    is_curtain[curtain_179]=True
    is_curtains[curtain_179]=True
    is_curtain[curtain_180]=True
    is_curtains[curtain_180]=True
    is_curtain[curtain_181]=True
    is_curtains[curtain_181]=True
    is_pillow[pillow_182]=True
    is_pillow[pillow_183]=True
    is_photoframe[photoframe_185]=True
    is_dining_room[dining_room_201]=True
    is_kitchen[dining_room_201]=True
    is_floor[floor_202]=True
    is_floor[floor_203]=True
    is_floor[floor_204]=True
    is_floor[floor_205]=True
    is_floor[floor_206]=True
    is_floor[floor_207]=True
    is_floor[floor_208]=True
    is_wall[wall_209]=True
    is_wall[wall_210]=True
    is_wall[wall_211]=True
    is_wall[wall_212]=True
    is_wall[wall_213]=True
    is_wall[wall_214]=True
    is_wall[wall_215]=True
    is_ceiling[ceiling_216]=True
    is_ceiling[ceiling_217]=True
    is_ceiling[ceiling_218]=True
    is_ceiling[ceiling_219]=True
    is_ceiling[ceiling_220]=True
    is_ceiling[ceiling_221]=True
    is_door[door_222]=True
    is_ceilinglamp[ceilinglamp_223]=True
    is_ceilinglamp[ceilinglamp_224]=True
    is_tvstand[tvstand_225]=True
    is_coffee_table[table_226]=True
    is_kitchen_table[table_226]=True
    is_table[table_226]=True
    is_diningtable[table_226]=True
    is_bench[bench_227]=True
    is_bench[bench_228]=True
    is_cupboard[cupboard_229]=True
    is_kitchen_cabinets[cupboard_229]=True
    is_kitchen_counter[kitchen_counter_230]=True
    is_sink[sink_231]=True
    is_faucet[faucet_232]=True
    is_bookshelf[bookshelf_233]=True
    is_wallshelf[wallshelf_234]=True
    is_wallshelf[wallshelf_235]=True
    is_rug[mat_236]=True
    is_mat[mat_236]=True
    is_rug[mat_237]=True
    is_mat[mat_237]=True
    is_wallpictureframe[drawing_238]=True
    is_drawing[drawing_238]=True
    is_wallpictureframe[drawing_239]=True
    is_drawing[drawing_239]=True
    is_wallpictureframe[drawing_240]=True
    is_drawing[drawing_240]=True
    is_wallpictureframe[drawing_241]=True
    is_drawing[drawing_241]=True
    is_wallpictureframe[drawing_242]=True
    is_drawing[drawing_242]=True
    is_wallpictureframe[drawing_243]=True
    is_drawing[drawing_243]=True
    is_orchid[orchid_244]=True
    is_light_switch[light_245]=True
    is_lightswitch[light_245]=True
    is_light[light_245]=True
    is_powersocket[powersocket_246]=True
    is_wall_phone[phone_247]=True
    is_phone[phone_247]=True
    is_cellphone[phone_247]=True
    is_television[television_248]=True
    is_tv[television_248]=True
    is_walltv[television_248]=True
    is_wall_clock[wall_clock_249]=True
    is_clock[wall_clock_249]=True
    is_photoframe[photoframe_285]=True
    is_stovefan[stovefan_288]=True
    is_freezer[fridge_289]=True
    is_fridge[fridge_289]=True
    is_coffeemaker[coffe_maker_290]=True
    is_coffe_maker[coffe_maker_290]=True
    is_toaster[toaster_292]=True
    is_stove[oven_295]=True
    is_oven[oven_295]=True
    is_tray[tray_296]=True
    is_oventray[tray_296]=True
    is_microwave[microwave_297]=True
    is_livingroom[home_office_319]=True
    is_home_office[home_office_319]=True
    is_floor[floor_320]=True
    is_floor[floor_321]=True
    is_floor[floor_322]=True
    is_floor[floor_323]=True
    is_floor[floor_324]=True
    is_floor[floor_325]=True
    is_floor[floor_326]=True
    is_floor[floor_327]=True
    is_floor[floor_328]=True
    is_wall[wall_329]=True
    is_wall[wall_330]=True
    is_wall[wall_331]=True
    is_wall[wall_332]=True
    is_wall[wall_333]=True
    is_wall[wall_334]=True
    is_wall[wall_335]=True
    is_wall[wall_336]=True
    is_ceiling[ceiling_337]=True
    is_ceiling[ceiling_338]=True
    is_ceiling[ceiling_339]=True
    is_ceiling[ceiling_340]=True
    is_ceiling[ceiling_341]=True
    is_ceiling[ceiling_342]=True
    is_ceiling[ceiling_343]=True
    is_ceiling[ceiling_344]=True
    is_ceiling[ceiling_345]=True
    is_doorjamb[doorjamb_346]=True
    is_doorjamb[doorjamb_347]=True
    is_window[window_348]=True
    is_ceilinglamp[ceilinglamp_349]=True
    is_walllamp[walllamp_350]=True
    is_walllamp[walllamp_351]=True
    is_couch[couch_352]=True
    is_sofa[couch_352]=True
    is_tvstand[tvstand_353]=True
    is_bookshelf[bookshelf_354]=True
    is_coffee_table[table_355]=True
    is_kitchen_table[table_355]=True
    is_table[table_355]=True
    is_diningtable[table_355]=True
    is_chair[chair_356]=True
    is_desk[desk_357]=True
    is_cpu_table[desk_357]=True
    is_closet[dresser_358]=True
    is_dresser[dresser_358]=True
    is_coatrack[hanger_359]=True
    is_hanger[hanger_359]=True
    is_coatrack[hanger_361]=True
    is_hanger[hanger_361]=True
    is_coatrack[hanger_363]=True
    is_hanger[hanger_363]=True
    is_coatrack[hanger_365]=True
    is_hanger[hanger_365]=True
    is_coatrack[hanger_367]=True
    is_hanger[hanger_367]=True
    is_coatrack[hanger_369]=True
    is_hanger[hanger_369]=True
    is_coatrack[hanger_372]=True
    is_hanger[hanger_372]=True
    is_coatrack[hanger_374]=True
    is_hanger[hanger_374]=True
    is_coatrack[hanger_375]=True
    is_hanger[hanger_375]=True
    is_coatrack[hanger_376]=True
    is_hanger[hanger_376]=True
    is_closetdrawer[closetdrawer_377]=True
    is_closetdrawer[closetdrawer_380]=True
    is_closetdrawer[closetdrawer_382]=True
    is_closetdrawer[closetdrawer_384]=True
    is_closetdrawer[closetdrawer_388]=True
    is_closetdrawer[closetdrawer_392]=True
    is_closetdrawer[closetdrawer_394]=True
    is_filing_cabinet[filing_cabinet_399]=True
    is_cabinet[filing_cabinet_399]=True
    is_wallpictureframe[drawing_400]=True
    is_drawing[drawing_400]=True
    is_rug[mat_401]=True
    is_mat[mat_401]=True
    is_wallpictureframe[drawing_402]=True
    is_drawing[drawing_402]=True
    is_wallpictureframe[drawing_403]=True
    is_drawing[drawing_403]=True
    is_wallpictureframe[drawing_404]=True
    is_drawing[drawing_404]=True
    is_pillow[pillow_405]=True
    is_pillow[pillow_406]=True
    is_curtain[curtain_407]=True
    is_curtains[curtain_407]=True
    is_curtain[curtain_408]=True
    is_curtains[curtain_408]=True
    is_curtain[curtain_409]=True
    is_curtains[curtain_409]=True
    is_television[television_410]=True
    is_tv[television_410]=True
    is_walltv[television_410]=True
    is_light_switch[light_411]=True
    is_lightswitch[light_411]=True
    is_light[light_411]=True
    is_powersocket[powersocket_412]=True
    is_mouse[mouse_413]=True
    is_mouse_mat[mousepad_414]=True
    is_mousemat[mousepad_414]=True
    is_mousepad[mousepad_414]=True
    is_keyboard[keyboard_415]=True
    is_cpuscreen[cpuscreen_416]=True
    is_cpu_case[computer_417]=True
    is_pc[computer_417]=True
    is_computer[computer_417]=True
    is_photoframe[photoframe_430]=True
    is_plate[plate_1000]=True
    is_dishwasher[dishwasher_1001]=True
    is_coffee_filter[coffee_filter_2000]=True
    is_pen[pencil_2001]=True
    is_pencil[pencil_2001]=True
    is_hairbrush[hairbrush_2002]=True
    is_wallpictureframe[drawing_2003]=True
    is_drawing[drawing_2003]=True
    is_chair[chair_2004]=True
    is_napkin[napkin_2005]=True
    is_cloth_napkin[napkin_2005]=True
    is_papertowel[napkin_2005]=True
    #categories_end

    #states
    is_on[ceilinglamp_26]=True
    is_on[walllamp_27]=True
    is_on[walllamp_28]=True
    is_on[walllamp_29]=True
    is_on[shower_36]=True
    is_on[ceilinglamp_96]=True
    is_on[tablelamp_97]=True
    is_on[tablelamp_98]=True
    is_on[ceilinglamp_223]=True
    is_on[ceilinglamp_224]=True
    is_on[fridge_289]=True
    is_on[oven_295]=True
    is_on[microwave_297]=True
    is_on[ceilinglamp_349]=True
    is_on[walllamp_350]=True
    is_on[walllamp_351]=True
    is_off[iron_2089]=True
    is_off[washing_machine_2007]=True
    is_off[remote_control_2052]=True
    is_off[cd_player_2060]=True
    is_off[dvd_player_2061]=True
    is_off[stove_2065]=True
    is_off[vacuum_cleaner_2070]=True
    is_off[phone_2077]=True
    is_off[toilet_37]=True
    is_off[faucet_43]=True
    is_off[light_64]=True
    is_off[light_169]=True
    is_off[computer_170]=True
    is_off[faucet_232]=True
    is_off[light_245]=True
    is_off[phone_247]=True
    is_off[television_248]=True
    is_off[wall_clock_249]=True
    is_off[coffe_maker_290]=True
    is_off[toaster_292]=True
    is_off[television_410]=True
    is_off[light_411]=True
    is_off[computer_417]=True
    is_off[dishwasher_1001]=True
    open[basket_for_clothes_2006]=True
    open[curtain_24]=True
    open[bathroom_counter_41]=True
    open[door_44]=True
    open[doorjamb_45]=True
    open[trashcan_99]=True
    open[nightstand_102]=True
    open[doorjamb_165]=True
    open[curtain_179]=True
    open[curtain_180]=True
    open[curtain_181]=True
    open[door_222]=True
    open[cupboard_229]=True
    open[doorjamb_346]=True
    open[doorjamb_347]=True
    open[curtain_407]=True
    closed[washing_machine_2007]=True
    closed[cd_player_2060]=True
    closed[dvd_player_2061]=True
    closed[stove_2065]=True
    closed[book_2066]=True
    closed[book_2067]=True
    closed[pot_2069]=True
    closed[curtain_23]=True
    closed[curtain_25]=True
    closed[toilet_37]=True
    closed[curtain_39]=True
    closed[bathroom_cabinet_40]=True
    closed[window_63]=True
    closed[light_64]=True
    closed[window_86]=True
    closed[nightstand_100]=True
    closed[bookshelf_101]=True
    closed[desk_104]=True
    closed[dresser_108]=True
    closed[dresser_123]=True
    closed[light_169]=True
    closed[kitchen_counter_230]=True
    closed[bookshelf_233]=True
    closed[light_245]=True
    closed[fridge_289]=True
    closed[coffe_maker_290]=True
    closed[oven_295]=True
    closed[microwave_297]=True
    closed[window_348]=True
    closed[bookshelf_354]=True
    closed[desk_357]=True
    closed[dresser_358]=True
    closed[filing_cabinet_399]=True
    closed[curtain_408]=True
    closed[curtain_409]=True
    closed[light_411]=True
    closed[dishwasher_1001]=True
    dirty[clothes_pants_2085]=True
    dirty[clothes_shirt_2086]=True
    dirty[clothes_socks_2087]=True
    dirty[clothes_skirt_2088]=True
    dirty[food_vegetable_2041]=True
    dirty[clothes_dress_2044]=True
    dirty[clothes_jacket_2047]=True
    dirty[clothes_scarf_2048]=True
    dirty[clothes_underwear_2049]=True
    dirty[bowl_2071]=True
    dirty[bowl_2072]=True
    dirty[floor_2]=True
    dirty[floor_4]=True
    dirty[floor_5]=True
    dirty[floor_7]=True
    dirty[floor_8]=True
    dirty[wall_9]=True
    dirty[wall_11]=True
    dirty[wall_12]=True
    dirty[wall_13]=True
    dirty[ceiling_19]=True
    dirty[ceiling_21]=True
    dirty[curtain_39]=True
    dirty[sink_42]=True
    dirty[window_63]=True
    dirty[floor_70]=True
    dirty[floor_71]=True
    dirty[floor_72]=True
    dirty[floor_73]=True
    dirty[floor_74]=True
    dirty[floor_77]=True
    dirty[wall_79]=True
    dirty[wall_80]=True
    dirty[wall_83]=True
    dirty[wall_84]=True
    dirty[wall_85]=True
    dirty[window_86]=True
    dirty[ceiling_88]=True
    dirty[ceiling_89]=True
    dirty[ceiling_92]=True
    dirty[ceiling_95]=True
    dirty[mousepad_167]=True
    dirty[floor_202]=True
    dirty[floor_205]=True
    dirty[floor_208]=True
    dirty[wall_209]=True
    dirty[wall_211]=True
    dirty[wall_212]=True
    dirty[ceiling_216]=True
    dirty[ceiling_217]=True
    dirty[ceiling_220]=True
    dirty[ceiling_221]=True
    dirty[table_226]=True
    dirty[sink_231]=True
    dirty[bookshelf_233]=True
    dirty[mat_236]=True
    dirty[floor_323]=True
    dirty[floor_328]=True
    dirty[wall_329]=True
    dirty[wall_330]=True
    dirty[wall_336]=True
    dirty[ceiling_339]=True
    dirty[ceiling_340]=True
    dirty[ceiling_343]=True
    dirty[ceiling_344]=True
    dirty[window_348]=True
    dirty[mat_401]=True
    dirty[pillow_405]=True
    dirty[curtain_409]=True
    dirty[plate_1000]=True
    clean[iron_2089]=True
    clean[washing_machine_2007]=True
    clean[food_steak_2008]=True
    clean[food_apple_2009]=True
    clean[food_bacon_2010]=True
    clean[food_banana_2011]=True
    clean[food_bread_2012]=True
    clean[food_cake_2013]=True
    clean[food_carrot_2014]=True
    clean[food_cereal_2015]=True
    clean[food_cheese_2016]=True
    clean[food_chicken_2017]=True
    clean[food_dessert_2018]=True
    clean[food_donut_2019]=True
    clean[food_egg_2020]=True
    clean[food_fish_2021]=True
    clean[food_food_2022]=True
    clean[food_fruit_2023]=True
    clean[food_hamburger_2024]=True
    clean[food_ice_cream_2025]=True
    clean[food_jam_2026]=True
    clean[food_kiwi_2027]=True
    clean[food_lemon_2028]=True
    clean[food_noodles_2029]=True
    clean[food_oatmeal_2030]=True
    clean[food_orange_2031]=True
    clean[food_onion_2032]=True
    clean[food_peanut_butter_2033]=True
    clean[food_pizza_2034]=True
    clean[food_potato_2035]=True
    clean[food_rice_2036]=True
    clean[food_salt_2037]=True
    clean[food_snack_2038]=True
    clean[food_sugar_2039]=True
    clean[food_turkey_2040]=True
    clean[dry_pasta_2042]=True
    clean[clothes_hat_2045]=True
    clean[clothes_gloves_2046]=True
    clean[knife_2050]=True
    clean[cutting_board_2051]=True
    clean[soap_2053]=True
    clean[soap_2054]=True
    clean[towel_2056]=True
    clean[towel_2057]=True
    clean[towel_2058]=True
    clean[towel_2059]=True
    clean[vacuum_cleaner_2070]=True
    clean[phone_2077]=True
    clean[fryingpan_2083]=True
    clean[detergent_2084]=True
    clean[bathroom_1]=True
    clean[floor_3]=True
    clean[floor_6]=True
    clean[wall_10]=True
    clean[wall_14]=True
    clean[wall_15]=True
    clean[ceiling_16]=True
    clean[ceiling_17]=True
    clean[ceiling_18]=True
    clean[ceiling_20]=True
    clean[mat_22]=True
    clean[curtain_23]=True
    clean[curtain_24]=True
    clean[curtain_25]=True
    clean[ceilinglamp_26]=True
    clean[walllamp_27]=True
    clean[walllamp_28]=True
    clean[walllamp_29]=True
    clean[bathtub_30]=True
    clean[towel_rack_31]=True
    clean[towel_rack_32]=True
    clean[towel_rack_33]=True
    clean[towel_rack_34]=True
    clean[wallshelf_35]=True
    clean[shower_36]=True
    clean[toilet_37]=True
    clean[shower_38]=True
    clean[bathroom_cabinet_40]=True
    clean[bathroom_counter_41]=True
    clean[faucet_43]=True
    clean[door_44]=True
    clean[doorjamb_45]=True
    clean[light_64]=True
    clean[bedroom_67]=True
    clean[floor_68]=True
    clean[floor_69]=True
    clean[floor_75]=True
    clean[floor_76]=True
    clean[wall_78]=True
    clean[wall_81]=True
    clean[wall_82]=True
    clean[ceiling_87]=True
    clean[ceiling_90]=True
    clean[ceiling_91]=True
    clean[ceiling_93]=True
    clean[ceiling_94]=True
    clean[ceilinglamp_96]=True
    clean[tablelamp_97]=True
    clean[tablelamp_98]=True
    clean[trashcan_99]=True
    clean[nightstand_100]=True
    clean[bookshelf_101]=True
    clean[nightstand_102]=True
    clean[chair_103]=True
    clean[desk_104]=True
    clean[bed_105]=True
    clean[chair_106]=True
    clean[table_107]=True
    clean[dresser_108]=True
    clean[hanger_109]=True
    clean[hanger_110]=True
    clean[hanger_111]=True
    clean[hanger_112]=True
    clean[hanger_113]=True
    clean[hanger_114]=True
    clean[hanger_115]=True
    clean[closetdrawer_116]=True
    clean[closetdrawer_117]=True
    clean[closetdrawer_118]=True
    clean[closetdrawer_119]=True
    clean[closetdrawer_120]=True
    clean[closetdrawer_121]=True
    clean[closetdrawer_122]=True
    clean[dresser_123]=True
    clean[hanger_124]=True
    clean[hanger_126]=True
    clean[hanger_128]=True
    clean[hanger_130]=True
    clean[hanger_132]=True
    clean[hanger_134]=True
    clean[hanger_136]=True
    clean[hanger_138]=True
    clean[hanger_140]=True
    clean[hanger_141]=True
    clean[hanger_142]=True
    clean[closetdrawer_143]=True
    clean[closetdrawer_146]=True
    clean[closetdrawer_148]=True
    clean[closetdrawer_150]=True
    clean[closetdrawer_154]=True
    clean[closetdrawer_158]=True
    clean[closetdrawer_160]=True
    clean[doorjamb_165]=True
    clean[mouse_166]=True
    clean[keyboard_168]=True
    clean[light_169]=True
    clean[computer_170]=True
    clean[cpuscreen_171]=True
    clean[mat_173]=True
    clean[drawing_174]=True
    clean[drawing_175]=True
    clean[drawing_176]=True
    clean[orchid_178]=True
    clean[curtain_179]=True
    clean[curtain_180]=True
    clean[curtain_181]=True
    clean[pillow_182]=True
    clean[pillow_183]=True
    clean[photoframe_185]=True
    clean[dining_room_201]=True
    clean[floor_203]=True
    clean[floor_204]=True
    clean[floor_206]=True
    clean[floor_207]=True
    clean[wall_210]=True
    clean[wall_213]=True
    clean[wall_214]=True
    clean[wall_215]=True
    clean[ceiling_218]=True
    clean[ceiling_219]=True
    clean[door_222]=True
    clean[ceilinglamp_223]=True
    clean[ceilinglamp_224]=True
    clean[tvstand_225]=True
    clean[bench_227]=True
    clean[bench_228]=True
    clean[cupboard_229]=True
    clean[kitchen_counter_230]=True
    clean[faucet_232]=True
    clean[wallshelf_234]=True
    clean[wallshelf_235]=True
    clean[mat_237]=True
    clean[drawing_238]=True
    clean[drawing_239]=True
    clean[drawing_240]=True
    clean[drawing_241]=True
    clean[drawing_242]=True
    clean[drawing_243]=True
    clean[orchid_244]=True
    clean[light_245]=True
    clean[powersocket_246]=True
    clean[phone_247]=True
    clean[television_248]=True
    clean[wall_clock_249]=True
    clean[photoframe_285]=True
    clean[stovefan_288]=True
    clean[fridge_289]=True
    clean[coffe_maker_290]=True
    clean[toaster_292]=True
    clean[oven_295]=True
    clean[tray_296]=True
    clean[microwave_297]=True
    clean[home_office_319]=True
    clean[floor_320]=True
    clean[floor_321]=True
    clean[floor_322]=True
    clean[floor_324]=True
    clean[floor_325]=True
    clean[floor_326]=True
    clean[floor_327]=True
    clean[wall_331]=True
    clean[wall_332]=True
    clean[wall_333]=True
    clean[wall_334]=True
    clean[wall_335]=True
    clean[ceiling_337]=True
    clean[ceiling_338]=True
    clean[ceiling_341]=True
    clean[ceiling_342]=True
    clean[ceiling_345]=True
    clean[doorjamb_346]=True
    clean[doorjamb_347]=True
    clean[ceilinglamp_349]=True
    clean[walllamp_350]=True
    clean[walllamp_351]=True
    clean[couch_352]=True
    clean[tvstand_353]=True
    clean[bookshelf_354]=True
    clean[table_355]=True
    clean[chair_356]=True
    clean[desk_357]=True
    clean[dresser_358]=True
    clean[hanger_359]=True
    clean[hanger_361]=True
    clean[hanger_363]=True
    clean[hanger_365]=True
    clean[hanger_367]=True
    clean[hanger_369]=True
    clean[hanger_372]=True
    clean[hanger_374]=True
    clean[hanger_375]=True
    clean[hanger_376]=True
    clean[closetdrawer_377]=True
    clean[closetdrawer_380]=True
    clean[closetdrawer_382]=True
    clean[closetdrawer_384]=True
    clean[closetdrawer_388]=True
    clean[closetdrawer_392]=True
    clean[closetdrawer_394]=True
    clean[filing_cabinet_399]=True
    clean[drawing_400]=True
    clean[drawing_402]=True
    clean[drawing_403]=True
    clean[drawing_404]=True
    clean[pillow_406]=True
    clean[curtain_407]=True
    clean[curtain_408]=True
    clean[television_410]=True
    clean[light_411]=True
    clean[powersocket_412]=True
    clean[mouse_413]=True
    clean[mousepad_414]=True
    clean[keyboard_415]=True
    clean[cpuscreen_416]=True
    clean[computer_417]=True
    clean[photoframe_430]=True
    clean[dishwasher_1001]=True
    clean[coffee_filter_2000]=True
    clean[pencil_2001]=True
    clean[hairbrush_2002]=True
    clean[drawing_2003]=True
    clean[chair_2004]=True
    clean[napkin_2005]=True
    plugged[light_64]=True
    plugged[keyboard_168]=True
    plugged[light_169]=True
    plugged[computer_170]=True
    plugged[light_245]=True
    plugged[television_248]=True
    plugged[wall_clock_249]=True
    plugged[fridge_289]=True
    plugged[coffe_maker_290]=True
    plugged[toaster_292]=True
    plugged[oven_295]=True
    plugged[microwave_297]=True
    plugged[television_410]=True
    plugged[light_411]=True
    plugged[mouse_413]=True
    plugged[keyboard_415]=True
    plugged[computer_417]=True
    plugged[dishwasher_1001]=True
    unplugged[iron_2089]=True
    unplugged[washing_machine_2007]=True
    unplugged[cd_player_2060]=True
    unplugged[dvd_player_2061]=True
    unplugged[vacuum_cleaner_2070]=True
    unplugged[mouse_166]=True
    unplugged[phone_247]=True
    used[cupboard_229]=True
    is_room[bathroom_1]=True
    is_room[bedroom_67]=True
    is_room[dining_room_201]=True
    is_room[home_office_319]=True
    #states_end

    #char_states
    standing[char]=True
    sitting[char]=False
    lying[char]=False
    sleeping[char]=False
    has_a_free_hand[char]=True
    #char_states_end

    #char
    close_char[char,wall_211]=True
    close_char[char,cupboard_229]=True
    inside_char[char,dining_room_201]=True
    #char_end

    #properties
    surfaces[cutting_board_2051]=True
    surfaces[cd_player_2060]=True
    surfaces[dvd_player_2061]=True
    surfaces[stove_2065]=True
    surfaces[coffee_table_2068]=True
    surfaces[ironing_board_2074]=True
    surfaces[floor_2]=True
    surfaces[floor_3]=True
    surfaces[floor_4]=True
    surfaces[floor_5]=True
    surfaces[floor_6]=True
    surfaces[floor_7]=True
    surfaces[floor_8]=True
    surfaces[mat_22]=True
    surfaces[towel_rack_31]=True
    surfaces[towel_rack_32]=True
    surfaces[towel_rack_33]=True
    surfaces[towel_rack_34]=True
    surfaces[bathroom_cabinet_40]=True
    surfaces[bathroom_counter_41]=True
    surfaces[floor_68]=True
    surfaces[floor_69]=True
    surfaces[floor_70]=True
    surfaces[floor_71]=True
    surfaces[floor_72]=True
    surfaces[floor_73]=True
    surfaces[floor_74]=True
    surfaces[floor_75]=True
    surfaces[floor_76]=True
    surfaces[floor_77]=True
    surfaces[nightstand_100]=True
    surfaces[bookshelf_101]=True
    surfaces[nightstand_102]=True
    surfaces[chair_103]=True
    surfaces[desk_104]=True
    surfaces[bed_105]=True
    surfaces[chair_106]=True
    surfaces[table_107]=True
    surfaces[mousepad_167]=True
    surfaces[mat_173]=True
    surfaces[floor_202]=True
    surfaces[floor_203]=True
    surfaces[floor_204]=True
    surfaces[floor_205]=True
    surfaces[floor_206]=True
    surfaces[floor_207]=True
    surfaces[floor_208]=True
    surfaces[tvstand_225]=True
    surfaces[table_226]=True
    surfaces[bench_227]=True
    surfaces[bench_228]=True
    surfaces[kitchen_counter_230]=True
    surfaces[bookshelf_233]=True
    surfaces[mat_236]=True
    surfaces[mat_237]=True
    surfaces[tray_296]=True
    surfaces[floor_320]=True
    surfaces[floor_321]=True
    surfaces[floor_322]=True
    surfaces[floor_323]=True
    surfaces[floor_324]=True
    surfaces[floor_325]=True
    surfaces[floor_326]=True
    surfaces[floor_327]=True
    surfaces[floor_328]=True
    surfaces[couch_352]=True
    surfaces[tvstand_353]=True
    surfaces[bookshelf_354]=True
    surfaces[table_355]=True
    surfaces[chair_356]=True
    surfaces[desk_357]=True
    surfaces[filing_cabinet_399]=True
    surfaces[mat_401]=True
    surfaces[mousepad_414]=True
    surfaces[plate_1000]=True
    surfaces[chair_2004]=True
    grabbable[clothes_pants_2085]=True
    grabbable[clothes_shirt_2086]=True
    grabbable[clothes_socks_2087]=True
    grabbable[clothes_skirt_2088]=True
    grabbable[iron_2089]=True
    grabbable[basket_for_clothes_2006]=True
    grabbable[food_steak_2008]=True
    grabbable[food_apple_2009]=True
    grabbable[food_bacon_2010]=True
    grabbable[food_banana_2011]=True
    grabbable[food_bread_2012]=True
    grabbable[food_cake_2013]=True
    grabbable[food_carrot_2014]=True
    grabbable[food_cereal_2015]=True
    grabbable[food_cheese_2016]=True
    grabbable[food_chicken_2017]=True
    grabbable[food_dessert_2018]=True
    grabbable[food_donut_2019]=True
    grabbable[food_egg_2020]=True
    grabbable[food_fish_2021]=True
    grabbable[food_food_2022]=True
    grabbable[food_fruit_2023]=True
    grabbable[food_hamburger_2024]=True
    grabbable[food_ice_cream_2025]=True
    grabbable[food_jam_2026]=True
    grabbable[food_kiwi_2027]=True
    grabbable[food_lemon_2028]=True
    grabbable[food_noodles_2029]=True
    grabbable[food_oatmeal_2030]=True
    grabbable[food_orange_2031]=True
    grabbable[food_onion_2032]=True
    grabbable[food_peanut_butter_2033]=True
    grabbable[food_pizza_2034]=True
    grabbable[food_potato_2035]=True
    grabbable[food_rice_2036]=True
    grabbable[food_salt_2037]=True
    grabbable[food_snack_2038]=True
    grabbable[food_sugar_2039]=True
    grabbable[food_turkey_2040]=True
    grabbable[food_vegetable_2041]=True
    grabbable[dry_pasta_2042]=True
    grabbable[milk_2043]=True
    grabbable[clothes_dress_2044]=True
    grabbable[clothes_hat_2045]=True
    grabbable[clothes_gloves_2046]=True
    grabbable[clothes_jacket_2047]=True
    grabbable[clothes_scarf_2048]=True
    grabbable[clothes_underwear_2049]=True
    grabbable[knife_2050]=True
    grabbable[cutting_board_2051]=True
    grabbable[remote_control_2052]=True
    grabbable[soap_2053]=True
    grabbable[soap_2054]=True
    grabbable[cat_2055]=True
    grabbable[towel_2056]=True
    grabbable[towel_2057]=True
    grabbable[towel_2058]=True
    grabbable[towel_2059]=True
    grabbable[cd_player_2060]=True
    grabbable[dvd_player_2061]=True
    grabbable[headset_2062]=True
    grabbable[cup_2063]=True
    grabbable[cup_2064]=True
    grabbable[book_2066]=True
    grabbable[book_2067]=True
    grabbable[pot_2069]=True
    grabbable[vacuum_cleaner_2070]=True
    grabbable[bowl_2071]=True
    grabbable[bowl_2072]=True
    grabbable[cleaning_solution_2073]=True
    grabbable[cd_2075]=True
    grabbable[headset_2076]=True
    grabbable[phone_2077]=True
    grabbable[sauce_2078]=True
    grabbable[oil_2079]=True
    grabbable[fork_2080]=True
    grabbable[fork_2081]=True
    grabbable[spectacles_2082]=True
    grabbable[fryingpan_2083]=True
    grabbable[detergent_2084]=True
    grabbable[mat_22]=True
    grabbable[towel_rack_31]=True
    grabbable[towel_rack_32]=True
    grabbable[towel_rack_33]=True
    grabbable[towel_rack_34]=True
    grabbable[chair_103]=True
    grabbable[chair_106]=True
    grabbable[hanger_109]=True
    grabbable[hanger_110]=True
    grabbable[hanger_111]=True
    grabbable[hanger_112]=True
    grabbable[hanger_113]=True
    grabbable[hanger_114]=True
    grabbable[hanger_115]=True
    grabbable[hanger_124]=True
    grabbable[hanger_126]=True
    grabbable[hanger_128]=True
    grabbable[hanger_130]=True
    grabbable[hanger_132]=True
    grabbable[hanger_134]=True
    grabbable[hanger_136]=True
    grabbable[hanger_138]=True
    grabbable[hanger_140]=True
    grabbable[hanger_141]=True
    grabbable[hanger_142]=True
    grabbable[mouse_166]=True
    grabbable[keyboard_168]=True
    grabbable[mat_173]=True
    grabbable[drawing_174]=True
    grabbable[drawing_175]=True
    grabbable[drawing_176]=True
    grabbable[pillow_182]=True
    grabbable[pillow_183]=True
    grabbable[mat_236]=True
    grabbable[mat_237]=True
    grabbable[drawing_238]=True
    grabbable[drawing_239]=True
    grabbable[drawing_240]=True
    grabbable[drawing_241]=True
    grabbable[drawing_242]=True
    grabbable[drawing_243]=True
    grabbable[phone_247]=True
    grabbable[wall_clock_249]=True
    grabbable[tray_296]=True
    grabbable[chair_356]=True
    grabbable[hanger_359]=True
    grabbable[hanger_361]=True
    grabbable[hanger_363]=True
    grabbable[hanger_365]=True
    grabbable[hanger_367]=True
    grabbable[hanger_369]=True
    grabbable[hanger_372]=True
    grabbable[hanger_374]=True
    grabbable[hanger_375]=True
    grabbable[hanger_376]=True
    grabbable[drawing_400]=True
    grabbable[mat_401]=True
    grabbable[drawing_402]=True
    grabbable[drawing_403]=True
    grabbable[drawing_404]=True
    grabbable[pillow_405]=True
    grabbable[pillow_406]=True
    grabbable[mouse_413]=True
    grabbable[keyboard_415]=True
    grabbable[plate_1000]=True
    grabbable[coffee_filter_2000]=True
    grabbable[pencil_2001]=True
    grabbable[hairbrush_2002]=True
    grabbable[drawing_2003]=True
    grabbable[chair_2004]=True
    grabbable[napkin_2005]=True
    sittable[mat_22]=True
    sittable[bathtub_30]=True
    sittable[toilet_37]=True
    sittable[chair_103]=True
    sittable[bed_105]=True
    sittable[chair_106]=True
    sittable[mat_173]=True
    sittable[bench_227]=True
    sittable[bench_228]=True
    sittable[mat_236]=True
    sittable[mat_237]=True
    sittable[couch_352]=True
    sittable[chair_356]=True
    sittable[mat_401]=True
    sittable[chair_2004]=True
    lieable[mat_22]=True
    lieable[bathtub_30]=True
    lieable[bed_105]=True
    lieable[mat_173]=True
    lieable[bench_227]=True
    lieable[bench_228]=True
    lieable[mat_236]=True
    lieable[mat_237]=True
    lieable[couch_352]=True
    lieable[mat_401]=True
    hangable[clothes_pants_2085]=True
    hangable[clothes_shirt_2086]=True
    hangable[clothes_socks_2087]=True
    hangable[clothes_skirt_2088]=True
    hangable[clothes_dress_2044]=True
    hangable[clothes_hat_2045]=True
    hangable[clothes_gloves_2046]=True
    hangable[clothes_jacket_2047]=True
    hangable[clothes_scarf_2048]=True
    hangable[clothes_underwear_2049]=True
    hangable[hanger_109]=True
    hangable[hanger_110]=True
    hangable[hanger_111]=True
    hangable[hanger_112]=True
    hangable[hanger_113]=True
    hangable[hanger_114]=True
    hangable[hanger_115]=True
    hangable[hanger_124]=True
    hangable[hanger_126]=True
    hangable[hanger_128]=True
    hangable[hanger_130]=True
    hangable[hanger_132]=True
    hangable[hanger_134]=True
    hangable[hanger_136]=True
    hangable[hanger_138]=True
    hangable[hanger_140]=True
    hangable[hanger_141]=True
    hangable[hanger_142]=True
    hangable[hanger_359]=True
    hangable[hanger_361]=True
    hangable[hanger_363]=True
    hangable[hanger_365]=True
    hangable[hanger_367]=True
    hangable[hanger_369]=True
    hangable[hanger_372]=True
    hangable[hanger_374]=True
    hangable[hanger_375]=True
    hangable[hanger_376]=True
    drinkable[milk_2043]=True
    drinkable[oil_2079]=True
    eatable[food_steak_2008]=True
    eatable[food_apple_2009]=True
    eatable[food_bacon_2010]=True
    eatable[food_banana_2011]=True
    eatable[food_bread_2012]=True
    eatable[food_cake_2013]=True
    eatable[food_carrot_2014]=True
    eatable[food_cereal_2015]=True
    eatable[food_cheese_2016]=True
    eatable[food_chicken_2017]=True
    eatable[food_dessert_2018]=True
    eatable[food_egg_2020]=True
    eatable[food_fish_2021]=True
    eatable[food_food_2022]=True
    eatable[food_fruit_2023]=True
    eatable[food_hamburger_2024]=True
    eatable[food_jam_2026]=True
    eatable[food_kiwi_2027]=True
    eatable[food_lemon_2028]=True
    eatable[food_noodles_2029]=True
    eatable[food_oatmeal_2030]=True
    eatable[food_orange_2031]=True
    eatable[food_onion_2032]=True
    eatable[food_peanut_butter_2033]=True
    eatable[food_pizza_2034]=True
    eatable[food_potato_2035]=True
    eatable[food_rice_2036]=True
    eatable[food_salt_2037]=True
    eatable[food_snack_2038]=True
    eatable[food_sugar_2039]=True
    eatable[food_turkey_2040]=True
    eatable[food_vegetable_2041]=True
    recipient[washing_machine_2007]=True
    recipient[cup_2063]=True
    recipient[cup_2064]=True
    recipient[pot_2069]=True
    recipient[bowl_2071]=True
    recipient[bowl_2072]=True
    recipient[fryingpan_2083]=True
    recipient[sink_42]=True
    recipient[sink_231]=True
    recipient[coffe_maker_290]=True
    recipient[plate_1000]=True
    cuttable[food_steak_2008]=True
    cuttable[food_apple_2009]=True
    cuttable[food_bacon_2010]=True
    cuttable[food_banana_2011]=True
    cuttable[food_bread_2012]=True
    cuttable[food_cake_2013]=True
    cuttable[food_carrot_2014]=True
    cuttable[food_cheese_2016]=True
    cuttable[food_chicken_2017]=True
    cuttable[food_dessert_2018]=True
    cuttable[food_egg_2020]=True
    cuttable[food_fish_2021]=True
    cuttable[food_food_2022]=True
    cuttable[food_fruit_2023]=True
    cuttable[food_hamburger_2024]=True
    cuttable[food_kiwi_2027]=True
    cuttable[food_lemon_2028]=True
    cuttable[food_orange_2031]=True
    cuttable[food_onion_2032]=True
    cuttable[food_pizza_2034]=True
    cuttable[food_potato_2035]=True
    cuttable[food_turkey_2040]=True
    cuttable[food_vegetable_2041]=True
    cuttable[book_2066]=True
    cuttable[book_2067]=True
    cuttable[drawing_174]=True
    cuttable[drawing_175]=True
    cuttable[drawing_176]=True
    cuttable[drawing_238]=True
    cuttable[drawing_239]=True
    cuttable[drawing_240]=True
    cuttable[drawing_241]=True
    cuttable[drawing_242]=True
    cuttable[drawing_243]=True
    cuttable[drawing_400]=True
    cuttable[drawing_402]=True
    cuttable[drawing_403]=True
    cuttable[drawing_404]=True
    cuttable[drawing_2003]=True
    pourable[food_cereal_2015]=True
    pourable[food_rice_2036]=True
    pourable[food_salt_2037]=True
    pourable[food_sugar_2039]=True
    pourable[milk_2043]=True
    pourable[cup_2063]=True
    pourable[cup_2064]=True
    pourable[cleaning_solution_2073]=True
    pourable[sauce_2078]=True
    pourable[oil_2079]=True
    pourable[detergent_2084]=True
    can_open[basket_for_clothes_2006]=True
    can_open[washing_machine_2007]=True
    can_open[food_cereal_2015]=True
    can_open[food_jam_2026]=True
    can_open[milk_2043]=True
    can_open[cd_player_2060]=True
    can_open[dvd_player_2061]=True
    can_open[stove_2065]=True
    can_open[book_2066]=True
    can_open[book_2067]=True
    can_open[pot_2069]=True
    can_open[curtain_23]=True
    can_open[curtain_24]=True
    can_open[curtain_25]=True
    can_open[toilet_37]=True
    can_open[curtain_39]=True
    can_open[bathroom_cabinet_40]=True
    can_open[door_44]=True
    can_open[window_63]=True
    can_open[window_86]=True
    can_open[trashcan_99]=True
    can_open[nightstand_100]=True
    can_open[bookshelf_101]=True
    can_open[nightstand_102]=True
    can_open[dresser_108]=True
    can_open[dresser_123]=True
    can_open[curtain_179]=True
    can_open[curtain_180]=True
    can_open[curtain_181]=True
    can_open[door_222]=True
    can_open[cupboard_229]=True
    can_open[bookshelf_233]=True
    can_open[fridge_289]=True
    can_open[coffe_maker_290]=True
    can_open[oven_295]=True
    can_open[microwave_297]=True
    can_open[window_348]=True
    can_open[bookshelf_354]=True
    can_open[dresser_358]=True
    can_open[filing_cabinet_399]=True
    can_open[curtain_407]=True
    can_open[curtain_408]=True
    can_open[curtain_409]=True
    can_open[dishwasher_1001]=True
    has_switch[iron_2089]=True
    has_switch[washing_machine_2007]=True
    has_switch[remote_control_2052]=True
    has_switch[cd_player_2060]=True
    has_switch[dvd_player_2061]=True
    has_switch[stove_2065]=True
    has_switch[vacuum_cleaner_2070]=True
    has_switch[phone_2077]=True
    has_switch[faucet_43]=True
    has_switch[light_64]=True
    has_switch[tablelamp_97]=True
    has_switch[tablelamp_98]=True
    has_switch[light_169]=True
    has_switch[computer_170]=True
    has_switch[faucet_232]=True
    has_switch[light_245]=True
    has_switch[phone_247]=True
    has_switch[television_248]=True
    has_switch[wall_clock_249]=True
    has_switch[fridge_289]=True
    has_switch[coffe_maker_290]=True
    has_switch[toaster_292]=True
    has_switch[oven_295]=True
    has_switch[microwave_297]=True
    has_switch[television_410]=True
    has_switch[light_411]=True
    has_switch[computer_417]=True
    has_switch[dishwasher_1001]=True
    containers[basket_for_clothes_2006]=True
    containers[washing_machine_2007]=True
    containers[cd_player_2060]=True
    containers[stove_2065]=True
    containers[pot_2069]=True
    containers[fryingpan_2083]=True
    containers[toilet_37]=True
    containers[bathroom_cabinet_40]=True
    containers[sink_42]=True
    containers[trashcan_99]=True
    containers[nightstand_100]=True
    containers[bookshelf_101]=True
    containers[nightstand_102]=True
    containers[dresser_108]=True
    containers[dresser_123]=True
    containers[cupboard_229]=True
    containers[sink_231]=True
    containers[bookshelf_233]=True
    containers[fridge_289]=True
    containers[coffe_maker_290]=True
    containers[toaster_292]=True
    containers[oven_295]=True
    containers[microwave_297]=True
    containers[bookshelf_354]=True
    containers[dresser_358]=True
    containers[filing_cabinet_399]=True
    containers[dishwasher_1001]=True
    has_plug[iron_2089]=True
    has_plug[washing_machine_2007]=True
    has_plug[cd_player_2060]=True
    has_plug[dvd_player_2061]=True
    has_plug[vacuum_cleaner_2070]=True
    has_plug[phone_2077]=True
    has_plug[light_64]=True
    has_plug[mouse_166]=True
    has_plug[keyboard_168]=True
    has_plug[light_169]=True
    has_plug[light_245]=True
    has_plug[phone_247]=True
    has_plug[television_248]=True
    has_plug[wall_clock_249]=True
    has_plug[fridge_289]=True
    has_plug[coffe_maker_290]=True
    has_plug[toaster_292]=True
    has_plug[oven_295]=True
    has_plug[microwave_297]=True
    has_plug[television_410]=True
    has_plug[light_411]=True
    has_plug[mouse_413]=True
    has_plug[keyboard_415]=True
    readable[book_2066]=True
    readable[book_2067]=True
    lookable[computer_170]=True
    lookable[drawing_174]=True
    lookable[drawing_175]=True
    lookable[drawing_176]=True
    lookable[drawing_238]=True
    lookable[drawing_239]=True
    lookable[drawing_240]=True
    lookable[drawing_241]=True
    lookable[drawing_242]=True
    lookable[drawing_243]=True
    lookable[television_248]=True
    lookable[wall_clock_249]=True
    lookable[drawing_400]=True
    lookable[drawing_402]=True
    lookable[drawing_403]=True
    lookable[drawing_404]=True
    lookable[television_410]=True
    lookable[computer_417]=True
    lookable[drawing_2003]=True
    is_clothes[clothes_pants_2085]=True
    is_clothes[clothes_shirt_2086]=True
    is_clothes[clothes_socks_2087]=True
    is_clothes[clothes_skirt_2088]=True
    is_clothes[clothes_dress_2044]=True
    is_clothes[clothes_hat_2045]=True
    is_clothes[clothes_gloves_2046]=True
    is_clothes[clothes_jacket_2047]=True
    is_clothes[clothes_scarf_2048]=True
    is_clothes[clothes_underwear_2049]=True
    is_clothes[headset_2062]=True
    is_clothes[headset_2076]=True
    is_clothes[spectacles_2082]=True
    is_food[food_steak_2008]=True
    is_food[food_apple_2009]=True
    is_food[food_bacon_2010]=True
    is_food[food_banana_2011]=True
    is_food[food_bread_2012]=True
    is_food[food_cake_2013]=True
    is_food[food_carrot_2014]=True
    is_food[food_cereal_2015]=True
    is_food[food_cheese_2016]=True
    is_food[food_chicken_2017]=True
    is_food[food_dessert_2018]=True
    is_food[food_donut_2019]=True
    is_food[food_egg_2020]=True
    is_food[food_fish_2021]=True
    is_food[food_food_2022]=True
    is_food[food_fruit_2023]=True
    is_food[food_hamburger_2024]=True
    is_food[food_ice_cream_2025]=True
    is_food[food_jam_2026]=True
    is_food[food_kiwi_2027]=True
    is_food[food_lemon_2028]=True
    is_food[food_noodles_2029]=True
    is_food[food_oatmeal_2030]=True
    is_food[food_orange_2031]=True
    is_food[food_onion_2032]=True
    is_food[food_peanut_butter_2033]=True
    is_food[food_pizza_2034]=True
    is_food[food_potato_2035]=True
    is_food[food_rice_2036]=True
    is_food[food_salt_2037]=True
    is_food[food_snack_2038]=True
    is_food[food_sugar_2039]=True
    is_food[food_turkey_2040]=True
    is_food[food_vegetable_2041]=True
    cover_object[towel_2056]=True
    cover_object[towel_2057]=True
    cover_object[towel_2058]=True
    cover_object[towel_2059]=True
    cover_object[curtain_23]=True
    cover_object[curtain_24]=True
    cover_object[curtain_25]=True
    cover_object[curtain_39]=True
    cover_object[curtain_179]=True
    cover_object[curtain_180]=True
    cover_object[curtain_181]=True
    cover_object[curtain_407]=True
    cover_object[curtain_408]=True
    cover_object[curtain_409]=True
    cover_object[napkin_2005]=True
    has_paper[book_2066]=True
    has_paper[book_2067]=True
    has_paper[drawing_174]=True
    has_paper[drawing_175]=True
    has_paper[drawing_176]=True
    has_paper[drawing_238]=True
    has_paper[drawing_239]=True
    has_paper[drawing_240]=True
    has_paper[drawing_241]=True
    has_paper[drawing_242]=True
    has_paper[drawing_243]=True
    has_paper[drawing_400]=True
    has_paper[drawing_402]=True
    has_paper[drawing_403]=True
    has_paper[drawing_404]=True
    has_paper[coffee_filter_2000]=True
    has_paper[drawing_2003]=True
    has_paper[napkin_2005]=True
    movable[clothes_pants_2085]=True
    movable[clothes_shirt_2086]=True
    movable[clothes_socks_2087]=True
    movable[clothes_skirt_2088]=True
    movable[iron_2089]=True
    movable[basket_for_clothes_2006]=True
    movable[food_steak_2008]=True
    movable[food_apple_2009]=True
    movable[food_bacon_2010]=True
    movable[food_banana_2011]=True
    movable[food_bread_2012]=True
    movable[food_cake_2013]=True
    movable[food_carrot_2014]=True
    movable[food_cereal_2015]=True
    movable[food_cheese_2016]=True
    movable[food_chicken_2017]=True
    movable[food_dessert_2018]=True
    movable[food_donut_2019]=True
    movable[food_egg_2020]=True
    movable[food_fish_2021]=True
    movable[food_food_2022]=True
    movable[food_fruit_2023]=True
    movable[food_hamburger_2024]=True
    movable[food_ice_cream_2025]=True
    movable[food_jam_2026]=True
    movable[food_kiwi_2027]=True
    movable[food_lemon_2028]=True
    movable[food_noodles_2029]=True
    movable[food_oatmeal_2030]=True
    movable[food_orange_2031]=True
    movable[food_onion_2032]=True
    movable[food_peanut_butter_2033]=True
    movable[food_pizza_2034]=True
    movable[food_potato_2035]=True
    movable[food_rice_2036]=True
    movable[food_salt_2037]=True
    movable[food_snack_2038]=True
    movable[food_sugar_2039]=True
    movable[food_turkey_2040]=True
    movable[food_vegetable_2041]=True
    movable[dry_pasta_2042]=True
    movable[milk_2043]=True
    movable[clothes_dress_2044]=True
    movable[clothes_hat_2045]=True
    movable[clothes_gloves_2046]=True
    movable[clothes_jacket_2047]=True
    movable[clothes_scarf_2048]=True
    movable[clothes_underwear_2049]=True
    movable[knife_2050]=True
    movable[cutting_board_2051]=True
    movable[remote_control_2052]=True
    movable[soap_2053]=True
    movable[soap_2054]=True
    movable[cat_2055]=True
    movable[towel_2056]=True
    movable[towel_2057]=True
    movable[towel_2058]=True
    movable[towel_2059]=True
    movable[cd_player_2060]=True
    movable[dvd_player_2061]=True
    movable[headset_2062]=True
    movable[cup_2063]=True
    movable[cup_2064]=True
    movable[book_2066]=True
    movable[book_2067]=True
    movable[coffee_table_2068]=True
    movable[pot_2069]=True
    movable[vacuum_cleaner_2070]=True
    movable[bowl_2071]=True
    movable[bowl_2072]=True
    movable[cleaning_solution_2073]=True
    movable[ironing_board_2074]=True
    movable[cd_2075]=True
    movable[headset_2076]=True
    movable[phone_2077]=True
    movable[sauce_2078]=True
    movable[oil_2079]=True
    movable[fork_2080]=True
    movable[fork_2081]=True
    movable[spectacles_2082]=True
    movable[fryingpan_2083]=True
    movable[detergent_2084]=True
    movable[mat_22]=True
    movable[curtain_23]=True
    movable[curtain_24]=True
    movable[curtain_25]=True
    movable[towel_rack_31]=True
    movable[towel_rack_32]=True
    movable[towel_rack_33]=True
    movable[towel_rack_34]=True
    movable[curtain_39]=True
    movable[trashcan_99]=True
    movable[chair_103]=True
    movable[desk_104]=True
    movable[chair_106]=True
    movable[table_107]=True
    movable[hanger_109]=True
    movable[hanger_110]=True
    movable[hanger_111]=True
    movable[hanger_112]=True
    movable[hanger_113]=True
    movable[hanger_114]=True
    movable[hanger_115]=True
    movable[hanger_124]=True
    movable[hanger_126]=True
    movable[hanger_128]=True
    movable[hanger_130]=True
    movable[hanger_132]=True
    movable[hanger_134]=True
    movable[hanger_136]=True
    movable[hanger_138]=True
    movable[hanger_140]=True
    movable[hanger_141]=True
    movable[hanger_142]=True
    movable[mouse_166]=True
    movable[mousepad_167]=True
    movable[keyboard_168]=True
    movable[mat_173]=True
    movable[drawing_174]=True
    movable[drawing_175]=True
    movable[drawing_176]=True
    movable[curtain_179]=True
    movable[curtain_180]=True
    movable[curtain_181]=True
    movable[pillow_182]=True
    movable[pillow_183]=True
    movable[table_226]=True
    movable[bench_227]=True
    movable[bench_228]=True
    movable[mat_236]=True
    movable[mat_237]=True
    movable[drawing_238]=True
    movable[drawing_239]=True
    movable[drawing_240]=True
    movable[drawing_241]=True
    movable[drawing_242]=True
    movable[drawing_243]=True
    movable[phone_247]=True
    movable[wall_clock_249]=True
    movable[coffe_maker_290]=True
    movable[toaster_292]=True
    movable[tray_296]=True
    movable[couch_352]=True
    movable[table_355]=True
    movable[chair_356]=True
    movable[desk_357]=True
    movable[hanger_359]=True
    movable[hanger_361]=True
    movable[hanger_363]=True
    movable[hanger_365]=True
    movable[hanger_367]=True
    movable[hanger_369]=True
    movable[hanger_372]=True
    movable[hanger_374]=True
    movable[hanger_375]=True
    movable[hanger_376]=True
    movable[drawing_400]=True
    movable[mat_401]=True
    movable[drawing_402]=True
    movable[drawing_403]=True
    movable[drawing_404]=True
    movable[pillow_405]=True
    movable[pillow_406]=True
    movable[curtain_407]=True
    movable[curtain_408]=True
    movable[curtain_409]=True
    movable[mouse_413]=True
    movable[mousepad_414]=True
    movable[keyboard_415]=True
    movable[plate_1000]=True
    movable[coffee_filter_2000]=True
    movable[pencil_2001]=True
    movable[hairbrush_2002]=True
    movable[drawing_2003]=True
    movable[chair_2004]=True
    movable[napkin_2005]=True
    cream[food_cheese_2016]=True
    cream[food_ice_cream_2025]=True
    cream[food_jam_2026]=True
    cream[food_peanut_butter_2033]=True
    cream[soap_2053]=True
    cream[soap_2054]=True
    cream[sauce_2078]=True
    has_size[cup_2063]=True
    has_size[cup_2064]=True
    has_size[coffe_maker_290]=True
    #properties_end

    #relations
    on[iron_2089,ironing_board_2074]=True
    on[clothes_dress_2044,bed_105]=True
    on[clothes_hat_2045,table_107]=True
    on[clothes_gloves_2046,table_107]=True
    on[clothes_jacket_2047,couch_352]=True
    on[knife_2050,kitchen_counter_230]=True
    on[cutting_board_2051,kitchen_counter_230]=True
    on[remote_control_2052,couch_352]=True
    on[soap_2053,sink_42]=True
    on[soap_2054,sink_231]=True
    on[cat_2055,couch_352]=True
    on[towel_2056,towel_rack_31]=True
    on[towel_2057,towel_rack_32]=True
    on[towel_2058,towel_rack_33]=True
    on[towel_2059,towel_rack_34]=True
    on[cd_player_2060,tvstand_225]=True
    on[dvd_player_2061,tvstand_353]=True
    on[headset_2062,table_355]=True
    on[cup_2063,kitchen_counter_230]=True
    on[cup_2064,kitchen_counter_230]=True
    on[stove_2065,kitchen_counter_230]=True
    on[book_2066,bookshelf_354]=True
    on[book_2067,bookshelf_354]=True
    on[pot_2069,kitchen_counter_230]=True
    on[bowl_2071,table_226]=True
    on[bowl_2072,table_226]=True
    on[cleaning_solution_2073,sink_42]=True
    on[cd_2075,tvstand_225]=True
    on[headset_2076,desk_357]=True
    on[phone_2077,desk_357]=True
    on[oil_2079,kitchen_counter_230]=True
    on[fork_2080,table_226]=True
    on[fork_2081,table_226]=True
    on[spectacles_2082,table_355]=True
    on[fryingpan_2083,kitchen_counter_230]=True
    on[detergent_2084,sink_42]=True
    on[ceiling_16,wall_12]=True
    on[ceiling_18,wall_11]=True
    on[ceiling_19,wall_10]=True
    on[ceiling_21,wall_9]=True
    on[bathtub_30,floor_5]=True
    on[bathroom_cabinet_40,wall_12]=True
    on[faucet_43,bathroom_counter_41]=True
    on[door_44,floor_6]=True
    on[door_44,floor_77]=True
    on[doorjamb_45,floor_6]=True
    on[ceiling_87,wall_81]=True
    on[ceiling_89,wall_82]=True
    on[ceiling_93,wall_83]=True
    on[ceiling_95,wall_85]=True
    on[tablelamp_97,nightstand_100]=True
    on[tablelamp_98,nightstand_102]=True
    on[nightstand_100,floor_69]=True
    on[nightstand_100,mat_173]=True
    on[bookshelf_101,floor_72]=True
    on[nightstand_102,floor_71]=True
    on[nightstand_102,mat_173]=True
    on[desk_104,floor_75]=True
    on[bed_105,floor_70]=True
    on[bed_105,mat_173]=True
    on[table_107,floor_73]=True
    on[closetdrawer_116,closetdrawer_119]=True
    on[closetdrawer_117,closetdrawer_118]=True
    on[closetdrawer_118,closetdrawer_121]=True
    on[closetdrawer_119,closetdrawer_120]=True
    on[closetdrawer_120,closetdrawer_122]=True
    on[closetdrawer_143,closetdrawer_150]=True
    on[closetdrawer_146,closetdrawer_148]=True
    on[closetdrawer_148,closetdrawer_158]=True
    on[closetdrawer_150,closetdrawer_154]=True
    on[closetdrawer_154,closetdrawer_160]=True
    on[mouse_166,desk_104]=True
    on[mouse_166,mousepad_167]=True
    on[mousepad_167,desk_104]=True
    on[keyboard_168,desk_104]=True
    on[cpuscreen_171,desk_104]=True
    on[orchid_178,table_107]=True
    on[pillow_182,bed_105]=True
    on[pillow_183,bed_105]=True
    on[ceiling_216,wall_211]=True
    on[ceiling_218,wall_210]=True
    on[ceiling_219,wall_213]=True
    on[ceiling_221,wall_212]=True
    on[door_222,floor_76]=True
    on[door_222,floor_206]=True
    on[tvstand_225,floor_208]=True
    on[bench_227,floor_205]=True
    on[bench_228,floor_205]=True
    on[cupboard_229,wall_211]=True
    on[faucet_232,kitchen_counter_230]=True
    on[bookshelf_233,floor_207]=True
    on[wallshelf_234,wall_212]=True
    on[mat_236,table_226]=True
    on[drawing_241,wall_214]=True
    on[orchid_244,tvstand_225]=True
    on[television_248,tvstand_225]=True
    on[photoframe_285,tvstand_225]=True
    on[fridge_289,floor_202]=True
    on[fridge_289,floor_203]=True
    on[coffe_maker_290,kitchen_counter_230]=True
    on[toaster_292,kitchen_counter_230]=True
    on[microwave_297,kitchen_counter_230]=True
    on[ceiling_337,wall_332]=True
    on[ceiling_339,wall_333]=True
    on[ceiling_343,wall_330]=True
    on[ceiling_345,wall_334]=True
    on[couch_352,mat_401]=True
    on[tvstand_353,floor_324]=True
    on[bookshelf_354,floor_320]=True
    on[table_355,mat_401]=True
    on[desk_357,floor_326]=True
    on[closetdrawer_377,closetdrawer_384]=True
    on[closetdrawer_380,closetdrawer_382]=True
    on[closetdrawer_382,closetdrawer_392]=True
    on[closetdrawer_384,closetdrawer_388]=True
    on[closetdrawer_388,closetdrawer_394]=True
    on[filing_cabinet_399,floor_320]=True
    on[drawing_404,wall_332]=True
    on[curtain_409,couch_352]=True
    on[television_410,tvstand_353]=True
    on[mouse_413,desk_357]=True
    on[mouse_413,mousepad_414]=True
    on[mousepad_414,desk_357]=True
    on[keyboard_415,desk_357]=True
    on[cpuscreen_416,desk_357]=True
    on[plate_1000,sink_231]=True
    on[coffee_filter_2000,table_226]=True
    on[pencil_2001,desk_357]=True
    on[hairbrush_2002,couch_352]=True
    on[drawing_2003,table_226]=True
    on[chair_2004,floor_69]=True
    on[napkin_2005,kitchen_counter_230]=True
    inside[clothes_pants_2085,basket_for_clothes_2006]=True
    inside[clothes_pants_2085,bathroom_1]=True
    inside[clothes_shirt_2086,basket_for_clothes_2006]=True
    inside[clothes_shirt_2086,bathroom_1]=True
    inside[clothes_socks_2087,basket_for_clothes_2006]=True
    inside[clothes_socks_2087,bathroom_1]=True
    inside[clothes_skirt_2088,basket_for_clothes_2006]=True
    inside[clothes_skirt_2088,bathroom_1]=True
    inside[iron_2089,bathroom_1]=True
    inside[basket_for_clothes_2006,bathroom_1]=True
    inside[washing_machine_2007,bathroom_1]=True
    inside[food_steak_2008,dining_room_201]=True
    inside[food_steak_2008,fridge_289]=True
    inside[food_apple_2009,dining_room_201]=True
    inside[food_apple_2009,fridge_289]=True
    inside[food_bacon_2010,dining_room_201]=True
    inside[food_bacon_2010,fridge_289]=True
    inside[food_banana_2011,dining_room_201]=True
    inside[food_banana_2011,fridge_289]=True
    inside[food_bread_2012,dining_room_201]=True
    inside[food_bread_2012,fridge_289]=True
    inside[food_cake_2013,dining_room_201]=True
    inside[food_cake_2013,fridge_289]=True
    inside[food_carrot_2014,dining_room_201]=True
    inside[food_carrot_2014,fridge_289]=True
    inside[food_cereal_2015,dining_room_201]=True
    inside[food_cereal_2015,fridge_289]=True
    inside[food_cheese_2016,dining_room_201]=True
    inside[food_cheese_2016,fridge_289]=True
    inside[food_chicken_2017,dining_room_201]=True
    inside[food_chicken_2017,fridge_289]=True
    inside[food_dessert_2018,dining_room_201]=True
    inside[food_dessert_2018,fridge_289]=True
    inside[food_donut_2019,dining_room_201]=True
    inside[food_donut_2019,fridge_289]=True
    inside[food_egg_2020,dining_room_201]=True
    inside[food_egg_2020,fridge_289]=True
    inside[food_fish_2021,dining_room_201]=True
    inside[food_fish_2021,fridge_289]=True
    inside[food_food_2022,dining_room_201]=True
    inside[food_food_2022,fridge_289]=True
    inside[food_fruit_2023,dining_room_201]=True
    inside[food_fruit_2023,fridge_289]=True
    inside[food_hamburger_2024,dining_room_201]=True
    inside[food_hamburger_2024,fridge_289]=True
    inside[food_ice_cream_2025,dining_room_201]=True
    inside[food_ice_cream_2025,fridge_289]=True
    inside[food_jam_2026,dining_room_201]=True
    inside[food_jam_2026,fridge_289]=True
    inside[food_kiwi_2027,dining_room_201]=True
    inside[food_kiwi_2027,fridge_289]=True
    inside[food_lemon_2028,dining_room_201]=True
    inside[food_lemon_2028,fridge_289]=True
    inside[food_noodles_2029,dining_room_201]=True
    inside[food_noodles_2029,fridge_289]=True
    inside[food_oatmeal_2030,dining_room_201]=True
    inside[food_oatmeal_2030,fridge_289]=True
    inside[food_orange_2031,dining_room_201]=True
    inside[food_orange_2031,fridge_289]=True
    inside[food_onion_2032,dining_room_201]=True
    inside[food_onion_2032,fridge_289]=True
    inside[food_peanut_butter_2033,dining_room_201]=True
    inside[food_peanut_butter_2033,fridge_289]=True
    inside[food_pizza_2034,dining_room_201]=True
    inside[food_pizza_2034,fridge_289]=True
    inside[food_potato_2035,dining_room_201]=True
    inside[food_potato_2035,fridge_289]=True
    inside[food_rice_2036,dining_room_201]=True
    inside[food_rice_2036,fridge_289]=True
    inside[food_salt_2037,dining_room_201]=True
    inside[food_salt_2037,fridge_289]=True
    inside[food_snack_2038,dining_room_201]=True
    inside[food_snack_2038,fridge_289]=True
    inside[food_sugar_2039,dining_room_201]=True
    inside[food_sugar_2039,fridge_289]=True
    inside[food_turkey_2040,dining_room_201]=True
    inside[food_turkey_2040,fridge_289]=True
    inside[food_vegetable_2041,dining_room_201]=True
    inside[food_vegetable_2041,fridge_289]=True
    inside[dry_pasta_2042,dining_room_201]=True
    inside[dry_pasta_2042,fridge_289]=True
    inside[milk_2043,dining_room_201]=True
    inside[milk_2043,fridge_289]=True
    inside[clothes_dress_2044,bedroom_67]=True
    inside[clothes_hat_2045,bedroom_67]=True
    inside[clothes_gloves_2046,bedroom_67]=True
    inside[clothes_jacket_2047,home_office_319]=True
    inside[clothes_scarf_2048,bedroom_67]=True
    inside[clothes_scarf_2048,bed_105]=True
    inside[clothes_underwear_2049,bedroom_67]=True
    inside[clothes_underwear_2049,bed_105]=True
    inside[knife_2050,dining_room_201]=True
    inside[cutting_board_2051,dining_room_201]=True
    inside[remote_control_2052,home_office_319]=True
    inside[soap_2053,bathroom_1]=True
    inside[soap_2054,dining_room_201]=True
    inside[cat_2055,home_office_319]=True
    inside[towel_2056,bathroom_1]=True
    inside[towel_2057,bathroom_1]=True
    inside[towel_2058,bathroom_1]=True
    inside[towel_2059,bathroom_1]=True
    inside[cd_player_2060,dining_room_201]=True
    inside[dvd_player_2061,home_office_319]=True
    inside[headset_2062,home_office_319]=True
    inside[cup_2063,dining_room_201]=True
    inside[cup_2064,dining_room_201]=True
    inside[stove_2065,dining_room_201]=True
    inside[book_2066,home_office_319]=True
    inside[book_2067,home_office_319]=True
    inside[coffee_table_2068,home_office_319]=True
    inside[pot_2069,dining_room_201]=True
    inside[vacuum_cleaner_2070,home_office_319]=True
    inside[bowl_2071,dining_room_201]=True
    inside[bowl_2072,dining_room_201]=True
    inside[cleaning_solution_2073,bathroom_1]=True
    inside[ironing_board_2074,bathroom_1]=True
    inside[cd_2075,dining_room_201]=True
    inside[headset_2076,home_office_319]=True
    inside[phone_2077,home_office_319]=True
    inside[sauce_2078,dining_room_201]=True
    inside[sauce_2078,fridge_289]=True
    inside[oil_2079,dining_room_201]=True
    inside[fork_2080,dining_room_201]=True
    inside[fork_2081,dining_room_201]=True
    inside[spectacles_2082,home_office_319]=True
    inside[fryingpan_2083,dining_room_201]=True
    inside[detergent_2084,bathroom_1]=True
    inside[floor_2,bathroom_1]=True
    inside[floor_3,bathroom_1]=True
    inside[floor_4,bathroom_1]=True
    inside[floor_5,bathroom_1]=True
    inside[floor_6,bathroom_1]=True
    inside[floor_7,bathroom_1]=True
    inside[floor_8,bathroom_1]=True
    inside[wall_9,bathroom_1]=True
    inside[wall_10,bathroom_1]=True
    inside[wall_11,bathroom_1]=True
    inside[wall_12,bathroom_1]=True
    inside[wall_13,bathroom_1]=True
    inside[wall_14,bathroom_1]=True
    inside[wall_15,bathroom_1]=True
    inside[ceiling_16,bathroom_1]=True
    inside[ceiling_17,bathroom_1]=True
    inside[ceiling_18,bathroom_1]=True
    inside[ceiling_19,bathroom_1]=True
    inside[ceiling_20,bathroom_1]=True
    inside[ceiling_21,bathroom_1]=True
    inside[mat_22,bathroom_1]=True
    inside[curtain_23,bathroom_1]=True
    inside[curtain_23,curtain_24]=True
    inside[curtain_24,bathroom_1]=True
    inside[curtain_24,curtain_23]=True
    inside[curtain_25,bathroom_1]=True
    inside[ceilinglamp_26,bathroom_1]=True
    inside[walllamp_27,bathroom_1]=True
    inside[walllamp_28,bathroom_1]=True
    inside[walllamp_29,bathroom_1]=True
    inside[bathtub_30,bathroom_1]=True
    inside[towel_rack_31,bathroom_1]=True
    inside[towel_rack_32,bathroom_1]=True
    inside[towel_rack_33,bathroom_1]=True
    inside[towel_rack_34,bathroom_1]=True
    inside[wallshelf_35,bathroom_1]=True
    inside[shower_36,bathroom_1]=True
    inside[toilet_37,bathroom_1]=True
    inside[shower_38,bathroom_1]=True
    inside[curtain_39,bathroom_1]=True
    inside[curtain_39,shower_38]=True
    inside[bathroom_cabinet_40,bathroom_1]=True
    inside[bathroom_counter_41,bathroom_1]=True
    inside[sink_42,bathroom_1]=True
    inside[sink_42,bathroom_counter_41]=True
    inside[faucet_43,bathroom_1]=True
    inside[door_44,bathroom_1]=True
    inside[doorjamb_45,bathroom_1]=True
    inside[window_63,bathroom_1]=True
    inside[light_64,bathroom_1]=True
    inside[floor_68,bedroom_67]=True
    inside[floor_69,bedroom_67]=True
    inside[floor_70,bedroom_67]=True
    inside[floor_71,bedroom_67]=True
    inside[floor_72,bedroom_67]=True
    inside[floor_73,bedroom_67]=True
    inside[floor_74,bedroom_67]=True
    inside[floor_75,bedroom_67]=True
    inside[floor_76,bedroom_67]=True
    inside[floor_77,bedroom_67]=True
    inside[wall_78,bedroom_67]=True
    inside[wall_79,bedroom_67]=True
    inside[wall_80,bedroom_67]=True
    inside[wall_81,bedroom_67]=True
    inside[wall_82,bedroom_67]=True
    inside[wall_83,bedroom_67]=True
    inside[wall_84,bedroom_67]=True
    inside[wall_85,bedroom_67]=True
    inside[window_86,bedroom_67]=True
    inside[ceiling_87,bedroom_67]=True
    inside[ceiling_88,bedroom_67]=True
    inside[ceiling_89,bedroom_67]=True
    inside[ceiling_90,bedroom_67]=True
    inside[ceiling_91,bedroom_67]=True
    inside[ceiling_92,bedroom_67]=True
    inside[ceiling_93,bedroom_67]=True
    inside[ceiling_94,bedroom_67]=True
    inside[ceiling_95,bedroom_67]=True
    inside[ceilinglamp_96,bedroom_67]=True
    inside[tablelamp_97,bedroom_67]=True
    inside[tablelamp_98,bedroom_67]=True
    inside[trashcan_99,bedroom_67]=True
    inside[nightstand_100,bedroom_67]=True
    inside[bookshelf_101,bedroom_67]=True
    inside[nightstand_102,bedroom_67]=True
    inside[chair_103,bedroom_67]=True
    inside[desk_104,bedroom_67]=True
    inside[bed_105,bedroom_67]=True
    inside[chair_106,bedroom_67]=True
    inside[table_107,bedroom_67]=True
    inside[dresser_108,bedroom_67]=True
    inside[hanger_109,bedroom_67]=True
    inside[hanger_109,dresser_108]=True
    inside[hanger_110,bedroom_67]=True
    inside[hanger_110,dresser_108]=True
    inside[hanger_111,bedroom_67]=True
    inside[hanger_111,dresser_108]=True
    inside[hanger_112,bedroom_67]=True
    inside[hanger_112,dresser_108]=True
    inside[hanger_113,bedroom_67]=True
    inside[hanger_113,dresser_108]=True
    inside[hanger_114,bedroom_67]=True
    inside[hanger_114,dresser_108]=True
    inside[hanger_115,bedroom_67]=True
    inside[hanger_115,dresser_108]=True
    inside[closetdrawer_116,bedroom_67]=True
    inside[closetdrawer_116,dresser_108]=True
    inside[closetdrawer_117,bedroom_67]=True
    inside[closetdrawer_117,dresser_108]=True
    inside[closetdrawer_118,bedroom_67]=True
    inside[closetdrawer_118,dresser_108]=True
    inside[closetdrawer_119,bedroom_67]=True
    inside[closetdrawer_119,dresser_108]=True
    inside[closetdrawer_120,bedroom_67]=True
    inside[closetdrawer_120,dresser_108]=True
    inside[closetdrawer_121,bedroom_67]=True
    inside[closetdrawer_121,dresser_108]=True
    inside[closetdrawer_122,bedroom_67]=True
    inside[closetdrawer_122,dresser_108]=True
    inside[dresser_123,bedroom_67]=True
    inside[hanger_124,bedroom_67]=True
    inside[hanger_124,dresser_123]=True
    inside[hanger_126,bedroom_67]=True
    inside[hanger_126,dresser_123]=True
    inside[hanger_128,bedroom_67]=True
    inside[hanger_128,dresser_123]=True
    inside[hanger_130,bedroom_67]=True
    inside[hanger_130,dresser_123]=True
    inside[hanger_132,bedroom_67]=True
    inside[hanger_132,dresser_123]=True
    inside[hanger_134,bedroom_67]=True
    inside[hanger_134,dresser_123]=True
    inside[hanger_136,bedroom_67]=True
    inside[hanger_136,dresser_123]=True
    inside[hanger_138,bedroom_67]=True
    inside[hanger_138,dresser_123]=True
    inside[hanger_140,bedroom_67]=True
    inside[hanger_140,dresser_123]=True
    inside[hanger_141,bedroom_67]=True
    inside[hanger_141,dresser_123]=True
    inside[hanger_142,bedroom_67]=True
    inside[hanger_142,dresser_123]=True
    inside[closetdrawer_143,bedroom_67]=True
    inside[closetdrawer_143,dresser_123]=True
    inside[closetdrawer_146,bedroom_67]=True
    inside[closetdrawer_146,dresser_123]=True
    inside[closetdrawer_148,bedroom_67]=True
    inside[closetdrawer_148,dresser_123]=True
    inside[closetdrawer_150,bedroom_67]=True
    inside[closetdrawer_150,dresser_123]=True
    inside[closetdrawer_154,bedroom_67]=True
    inside[closetdrawer_154,dresser_123]=True
    inside[closetdrawer_158,bedroom_67]=True
    inside[closetdrawer_158,dresser_123]=True
    inside[closetdrawer_160,bedroom_67]=True
    inside[closetdrawer_160,dresser_123]=True
    inside[doorjamb_165,bedroom_67]=True
    inside[mouse_166,bedroom_67]=True
    inside[mousepad_167,bedroom_67]=True
    inside[keyboard_168,bedroom_67]=True
    inside[light_169,bedroom_67]=True
    inside[computer_170,bedroom_67]=True
    inside[cpuscreen_171,bedroom_67]=True
    inside[mat_173,bedroom_67]=True
    inside[drawing_174,bedroom_67]=True
    inside[drawing_175,bedroom_67]=True
    inside[drawing_176,bedroom_67]=True
    inside[orchid_178,bedroom_67]=True
    inside[curtain_179,bedroom_67]=True
    inside[curtain_179,curtain_180]=True
    inside[curtain_180,bedroom_67]=True
    inside[curtain_180,curtain_179]=True
    inside[curtain_181,bedroom_67]=True
    inside[pillow_182,bedroom_67]=True
    inside[pillow_183,bedroom_67]=True
    inside[photoframe_185,bedroom_67]=True
    inside[photoframe_185,bookshelf_101]=True
    inside[floor_202,dining_room_201]=True
    inside[floor_203,dining_room_201]=True
    inside[floor_204,dining_room_201]=True
    inside[floor_205,dining_room_201]=True
    inside[floor_206,dining_room_201]=True
    inside[floor_207,dining_room_201]=True
    inside[floor_208,dining_room_201]=True
    inside[wall_209,dining_room_201]=True
    inside[wall_210,dining_room_201]=True
    inside[wall_211,dining_room_201]=True
    inside[wall_212,dining_room_201]=True
    inside[wall_213,dining_room_201]=True
    inside[wall_214,dining_room_201]=True
    inside[wall_215,dining_room_201]=True
    inside[ceiling_216,dining_room_201]=True
    inside[ceiling_217,dining_room_201]=True
    inside[ceiling_218,dining_room_201]=True
    inside[ceiling_219,dining_room_201]=True
    inside[ceiling_220,dining_room_201]=True
    inside[ceiling_221,dining_room_201]=True
    inside[door_222,dining_room_201]=True
    inside[ceilinglamp_223,dining_room_201]=True
    inside[ceilinglamp_224,dining_room_201]=True
    inside[tvstand_225,dining_room_201]=True
    inside[table_226,dining_room_201]=True
    inside[bench_227,dining_room_201]=True
    inside[bench_228,dining_room_201]=True
    inside[cupboard_229,dining_room_201]=True
    inside[kitchen_counter_230,dining_room_201]=True
    inside[sink_231,dining_room_201]=True
    inside[sink_231,kitchen_counter_230]=True
    inside[faucet_232,dining_room_201]=True
    inside[bookshelf_233,dining_room_201]=True
    inside[wallshelf_234,dining_room_201]=True
    inside[wallshelf_235,dining_room_201]=True
    inside[mat_236,dining_room_201]=True
    inside[mat_237,dining_room_201]=True
    inside[drawing_238,dining_room_201]=True
    inside[drawing_239,dining_room_201]=True
    inside[drawing_240,dining_room_201]=True
    inside[drawing_241,dining_room_201]=True
    inside[drawing_242,dining_room_201]=True
    inside[drawing_243,dining_room_201]=True
    inside[orchid_244,dining_room_201]=True
    inside[light_245,dining_room_201]=True
    inside[powersocket_246,dining_room_201]=True
    inside[phone_247,dining_room_201]=True
    inside[television_248,dining_room_201]=True
    inside[wall_clock_249,dining_room_201]=True
    inside[photoframe_285,dining_room_201]=True
    inside[stovefan_288,dining_room_201]=True
    inside[fridge_289,dining_room_201]=True
    inside[coffe_maker_290,dining_room_201]=True
    inside[toaster_292,dining_room_201]=True
    inside[oven_295,dining_room_201]=True
    inside[tray_296,dining_room_201]=True
    inside[tray_296,oven_295]=True
    inside[microwave_297,dining_room_201]=True
    inside[floor_320,home_office_319]=True
    inside[floor_321,home_office_319]=True
    inside[floor_322,home_office_319]=True
    inside[floor_323,home_office_319]=True
    inside[floor_324,home_office_319]=True
    inside[floor_325,home_office_319]=True
    inside[floor_326,home_office_319]=True
    inside[floor_327,home_office_319]=True
    inside[floor_328,home_office_319]=True
    inside[wall_329,home_office_319]=True
    inside[wall_330,home_office_319]=True
    inside[wall_331,home_office_319]=True
    inside[wall_332,home_office_319]=True
    inside[wall_333,home_office_319]=True
    inside[wall_334,home_office_319]=True
    inside[wall_335,home_office_319]=True
    inside[wall_336,home_office_319]=True
    inside[ceiling_337,home_office_319]=True
    inside[ceiling_338,home_office_319]=True
    inside[ceiling_339,home_office_319]=True
    inside[ceiling_340,home_office_319]=True
    inside[ceiling_341,home_office_319]=True
    inside[ceiling_342,home_office_319]=True
    inside[ceiling_343,home_office_319]=True
    inside[ceiling_344,home_office_319]=True
    inside[ceiling_345,home_office_319]=True
    inside[doorjamb_346,home_office_319]=True
    inside[doorjamb_347,home_office_319]=True
    inside[window_348,home_office_319]=True
    inside[ceilinglamp_349,home_office_319]=True
    inside[walllamp_350,home_office_319]=True
    inside[walllamp_351,home_office_319]=True
    inside[couch_352,home_office_319]=True
    inside[tvstand_353,home_office_319]=True
    inside[bookshelf_354,home_office_319]=True
    inside[table_355,home_office_319]=True
    inside[table_355,couch_352]=True
    inside[chair_356,home_office_319]=True
    inside[desk_357,home_office_319]=True
    inside[dresser_358,home_office_319]=True
    inside[hanger_359,home_office_319]=True
    inside[hanger_359,dresser_358]=True
    inside[hanger_361,home_office_319]=True
    inside[hanger_361,dresser_358]=True
    inside[hanger_363,home_office_319]=True
    inside[hanger_363,dresser_358]=True
    inside[hanger_365,home_office_319]=True
    inside[hanger_365,dresser_358]=True
    inside[hanger_367,home_office_319]=True
    inside[hanger_367,dresser_358]=True
    inside[hanger_369,home_office_319]=True
    inside[hanger_369,dresser_358]=True
    inside[hanger_372,home_office_319]=True
    inside[hanger_372,dresser_358]=True
    inside[hanger_374,home_office_319]=True
    inside[hanger_374,dresser_358]=True
    inside[hanger_375,home_office_319]=True
    inside[hanger_375,dresser_358]=True
    inside[hanger_376,home_office_319]=True
    inside[hanger_376,dresser_358]=True
    inside[closetdrawer_377,home_office_319]=True
    inside[closetdrawer_377,dresser_358]=True
    inside[closetdrawer_380,home_office_319]=True
    inside[closetdrawer_380,dresser_358]=True
    inside[closetdrawer_382,home_office_319]=True
    inside[closetdrawer_382,dresser_358]=True
    inside[closetdrawer_384,home_office_319]=True
    inside[closetdrawer_384,dresser_358]=True
    inside[closetdrawer_388,home_office_319]=True
    inside[closetdrawer_388,dresser_358]=True
    inside[closetdrawer_392,home_office_319]=True
    inside[closetdrawer_392,dresser_358]=True
    inside[closetdrawer_394,home_office_319]=True
    inside[closetdrawer_394,dresser_358]=True
    inside[filing_cabinet_399,home_office_319]=True
    inside[drawing_400,home_office_319]=True
    inside[mat_401,home_office_319]=True
    inside[drawing_402,home_office_319]=True
    inside[drawing_403,home_office_319]=True
    inside[drawing_404,home_office_319]=True
    inside[pillow_405,home_office_319]=True
    inside[pillow_406,home_office_319]=True
    inside[pillow_406,couch_352]=True
    inside[curtain_407,home_office_319]=True
    inside[curtain_407,curtain_408]=True
    inside[curtain_408,home_office_319]=True
    inside[curtain_408,curtain_407]=True
    inside[curtain_409,home_office_319]=True
    inside[television_410,home_office_319]=True
    inside[light_411,home_office_319]=True
    inside[powersocket_412,home_office_319]=True
    inside[mouse_413,home_office_319]=True
    inside[mousepad_414,home_office_319]=True
    inside[keyboard_415,home_office_319]=True
    inside[cpuscreen_416,home_office_319]=True
    inside[computer_417,home_office_319]=True
    inside[photoframe_430,home_office_319]=True
    inside[photoframe_430,bookshelf_354]=True
    inside[plate_1000,dining_room_201]=True
    inside[dishwasher_1001,dining_room_201]=True
    inside[coffee_filter_2000,dining_room_201]=True
    inside[pencil_2001,home_office_319]=True
    inside[hairbrush_2002,home_office_319]=True
    inside[drawing_2003,dining_room_201]=True
    inside[chair_2004,bedroom_67]=True
    inside[napkin_2005,dining_room_201]=True
    between[door_44,bathroom_1]=True
    between[door_44,bedroom_67]=True
    between[door_222,bedroom_67]=True
    between[door_222,dining_room_201]=True
    between[doorjamb_346,dining_room_201]=True
    between[doorjamb_346,home_office_319]=True
    close[clothes_pants_2085,basket_for_clothes_2006]=True
    close[clothes_shirt_2086,basket_for_clothes_2006]=True
    close[clothes_socks_2087,basket_for_clothes_2006]=True
    close[clothes_skirt_2088,basket_for_clothes_2006]=True
    close[iron_2089,ironing_board_2074]=True
    close[basket_for_clothes_2006,clothes_pants_2085]=True
    close[basket_for_clothes_2006,clothes_shirt_2086]=True
    close[basket_for_clothes_2006,clothes_socks_2087]=True
    close[basket_for_clothes_2006,clothes_skirt_2088]=True
    close[basket_for_clothes_2006,mat_22]=True
    close[basket_for_clothes_2006,bathtub_30]=True
    close[basket_for_clothes_2006,towel_rack_31]=True
    close[basket_for_clothes_2006,towel_rack_32]=True
    close[basket_for_clothes_2006,towel_rack_33]=True
    close[basket_for_clothes_2006,towel_rack_34]=True
    close[basket_for_clothes_2006,shower_36]=True
    close[basket_for_clothes_2006,toilet_37]=True
    close[basket_for_clothes_2006,sink_42]=True
    close[basket_for_clothes_2006,faucet_43]=True
    close[washing_machine_2007,sink_42]=True
    close[food_steak_2008,fridge_289]=True
    close[food_apple_2009,fridge_289]=True
    close[food_bacon_2010,fridge_289]=True
    close[food_banana_2011,fridge_289]=True
    close[food_bread_2012,fridge_289]=True
    close[food_cake_2013,fridge_289]=True
    close[food_carrot_2014,fridge_289]=True
    close[food_cereal_2015,fridge_289]=True
    close[food_cheese_2016,fridge_289]=True
    close[food_chicken_2017,fridge_289]=True
    close[food_dessert_2018,fridge_289]=True
    close[food_donut_2019,fridge_289]=True
    close[food_egg_2020,fridge_289]=True
    close[food_fish_2021,fridge_289]=True
    close[food_food_2022,fridge_289]=True
    close[food_fruit_2023,fridge_289]=True
    close[food_hamburger_2024,fridge_289]=True
    close[food_ice_cream_2025,fridge_289]=True
    close[food_jam_2026,fridge_289]=True
    close[food_kiwi_2027,fridge_289]=True
    close[food_lemon_2028,fridge_289]=True
    close[food_noodles_2029,fridge_289]=True
    close[food_oatmeal_2030,fridge_289]=True
    close[food_orange_2031,fridge_289]=True
    close[food_onion_2032,fridge_289]=True
    close[food_peanut_butter_2033,fridge_289]=True
    close[food_pizza_2034,fridge_289]=True
    close[food_potato_2035,fridge_289]=True
    close[food_rice_2036,fridge_289]=True
    close[food_salt_2037,fridge_289]=True
    close[food_snack_2038,fridge_289]=True
    close[food_sugar_2039,fridge_289]=True
    close[food_turkey_2040,fridge_289]=True
    close[food_vegetable_2041,fridge_289]=True
    close[dry_pasta_2042,fridge_289]=True
    close[milk_2043,fridge_289]=True
    close[clothes_dress_2044,bed_105]=True
    close[clothes_hat_2045,table_107]=True
    close[clothes_gloves_2046,table_107]=True
    close[clothes_jacket_2047,couch_352]=True
    close[clothes_scarf_2048,bed_105]=True
    close[clothes_underwear_2049,bed_105]=True
    close[knife_2050,kitchen_counter_230]=True
    close[cutting_board_2051,kitchen_counter_230]=True
    close[remote_control_2052,couch_352]=True
    close[soap_2053,sink_42]=True
    close[soap_2054,sink_231]=True
    close[cat_2055,couch_352]=True
    close[towel_2056,towel_rack_31]=True
    close[towel_2057,towel_rack_32]=True
    close[towel_2058,towel_rack_33]=True
    close[towel_2059,towel_rack_34]=True
    close[cd_player_2060,tvstand_225]=True
    close[dvd_player_2061,tvstand_353]=True
    close[headset_2062,table_355]=True
    close[cup_2063,kitchen_counter_230]=True
    close[cup_2064,kitchen_counter_230]=True
    close[stove_2065,kitchen_counter_230]=True
    close[book_2066,bookshelf_354]=True
    close[book_2067,bookshelf_354]=True
    close[coffee_table_2068,home_office_319]=True
    close[pot_2069,kitchen_counter_230]=True
    close[vacuum_cleaner_2070,couch_352]=True
    close[bowl_2071,table_226]=True
    close[bowl_2072,table_226]=True
    close[cleaning_solution_2073,sink_42]=True
    close[ironing_board_2074,iron_2089]=True
    close[ironing_board_2074,bathroom_1]=True
    close[cd_2075,tvstand_225]=True
    close[headset_2076,desk_357]=True
    close[phone_2077,desk_357]=True
    close[sauce_2078,fridge_289]=True
    close[oil_2079,kitchen_counter_230]=True
    close[fork_2080,table_226]=True
    close[fork_2081,table_226]=True
    close[spectacles_2082,table_355]=True
    close[fryingpan_2083,kitchen_counter_230]=True
    close[detergent_2084,sink_42]=True
    close[bathroom_1,ironing_board_2074]=True
    close[floor_2,floor_3]=True
    close[floor_2,floor_4]=True
    close[floor_2,floor_6]=True
    close[floor_2,wall_9]=True
    close[floor_2,wall_12]=True
    close[floor_2,mat_22]=True
    close[floor_2,walllamp_28]=True
    close[floor_2,towel_rack_31]=True
    close[floor_2,towel_rack_32]=True
    close[floor_2,bathroom_counter_41]=True
    close[floor_2,sink_42]=True
    close[floor_2,faucet_43]=True
    close[floor_2,door_44]=True
    close[floor_2,light_64]=True
    close[floor_2,floor_72]=True
    close[floor_2,wall_79]=True
    close[floor_2,bookshelf_101]=True
    close[floor_2,drawing_176]=True
    close[floor_3,floor_2]=True
    close[floor_3,floor_4]=True
    close[floor_3,floor_6]=True
    close[floor_3,wall_9]=True
    close[floor_3,wall_12]=True
    close[floor_3,mat_22]=True
    close[floor_3,walllamp_28]=True
    close[floor_3,towel_rack_31]=True
    close[floor_3,towel_rack_32]=True
    close[floor_3,bathroom_counter_41]=True
    close[floor_3,sink_42]=True
    close[floor_3,faucet_43]=True
    close[floor_3,door_44]=True
    close[floor_3,light_64]=True
    close[floor_3,floor_72]=True
    close[floor_3,wall_79]=True
    close[floor_3,bookshelf_101]=True
    close[floor_3,drawing_176]=True
    close[floor_4,floor_2]=True
    close[floor_4,floor_3]=True
    close[floor_4,floor_5]=True
    close[floor_4,wall_9]=True
    close[floor_4,wall_12]=True
    close[floor_4,walllamp_27]=True
    close[floor_4,bathtub_30]=True
    close[floor_4,towel_rack_33]=True
    close[floor_4,towel_rack_34]=True
    close[floor_4,bathroom_counter_41]=True
    close[floor_4,sink_42]=True
    close[floor_4,faucet_43]=True
    close[floor_5,floor_4]=True
    close[floor_5,floor_6]=True
    close[floor_5,floor_8]=True
    close[floor_5,wall_9]=True
    close[floor_5,wall_10]=True
    close[floor_5,wall_13]=True
    close[floor_5,mat_22]=True
    close[floor_5,curtain_23]=True
    close[floor_5,curtain_24]=True
    close[floor_5,curtain_25]=True
    close[floor_5,bathtub_30]=True
    close[floor_5,towel_rack_33]=True
    close[floor_5,window_63]=True
    close[floor_6,floor_2]=True
    close[floor_6,floor_3]=True
    close[floor_6,floor_5]=True
    close[floor_6,floor_7]=True
    close[floor_6,wall_11]=True
    close[floor_6,wall_12]=True
    close[floor_6,wall_14]=True
    close[floor_6,mat_22]=True
    close[floor_6,towel_rack_32]=True
    close[floor_6,door_44]=True
    close[floor_6,doorjamb_45]=True
    close[floor_6,light_64]=True
    close[floor_6,floor_77]=True
    close[floor_6,wall_85]=True
    close[floor_6,fridge_289]=True
    close[floor_7,floor_6]=True
    close[floor_7,floor_8]=True
    close[floor_7,wall_10]=True
    close[floor_7,wall_11]=True
    close[floor_7,wall_15]=True
    close[floor_7,mat_22]=True
    close[floor_7,walllamp_29]=True
    close[floor_7,shower_36]=True
    close[floor_7,toilet_37]=True
    close[floor_7,door_44]=True
    close[floor_7,floor_202]=True
    close[floor_7,floor_203]=True
    close[floor_7,wall_211]=True
    close[floor_7,kitchen_counter_230]=True
    close[floor_7,sink_231]=True
    close[floor_7,faucet_232]=True
    close[floor_7,fridge_289]=True
    close[floor_7,toaster_292]=True
    close[floor_7,microwave_297]=True
    close[floor_8,floor_5]=True
    close[floor_8,floor_7]=True
    close[floor_8,wall_10]=True
    close[floor_8,wall_11]=True
    close[floor_8,walllamp_29]=True
    close[floor_8,bathtub_30]=True
    close[floor_8,shower_38]=True
    close[floor_8,curtain_39]=True
    close[wall_9,floor_2]=True
    close[wall_9,floor_3]=True
    close[wall_9,floor_4]=True
    close[wall_9,floor_5]=True
    close[wall_9,wall_12]=True
    close[wall_9,wall_13]=True
    close[wall_9,ceiling_16]=True
    close[wall_9,ceiling_20]=True
    close[wall_9,ceiling_21]=True
    close[wall_9,curtain_23]=True
    close[wall_9,curtain_24]=True
    close[wall_9,ceilinglamp_26]=True
    close[wall_9,walllamp_27]=True
    close[wall_9,bathtub_30]=True
    close[wall_9,towel_rack_33]=True
    close[wall_9,towel_rack_34]=True
    close[wall_9,wallshelf_35]=True
    close[wall_9,bathroom_cabinet_40]=True
    close[wall_9,bathroom_counter_41]=True
    close[wall_9,sink_42]=True
    close[wall_9,faucet_43]=True
    close[wall_9,window_63]=True
    close[wall_10,floor_5]=True
    close[wall_10,floor_7]=True
    close[wall_10,floor_8]=True
    close[wall_10,wall_11]=True
    close[wall_10,wall_13]=True
    close[wall_10,ceiling_18]=True
    close[wall_10,ceiling_19]=True
    close[wall_10,ceiling_20]=True
    close[wall_10,curtain_25]=True
    close[wall_10,ceilinglamp_26]=True
    close[wall_10,walllamp_29]=True
    close[wall_10,bathtub_30]=True
    close[wall_10,shower_38]=True
    close[wall_10,curtain_39]=True
    close[wall_10,window_63]=True
    close[wall_11,floor_6]=True
    close[wall_11,floor_7]=True
    close[wall_11,floor_8]=True
    close[wall_11,wall_10]=True
    close[wall_11,wall_14]=True
    close[wall_11,wall_15]=True
    close[wall_11,ceiling_17]=True
    close[wall_11,ceiling_18]=True
    close[wall_11,ceiling_19]=True
    close[wall_11,mat_22]=True
    close[wall_11,ceilinglamp_26]=True
    close[wall_11,walllamp_29]=True
    close[wall_11,shower_36]=True
    close[wall_11,toilet_37]=True
    close[wall_11,curtain_39]=True
    close[wall_11,door_44]=True
    close[wall_11,doorjamb_45]=True
    close[wall_11,floor_202]=True
    close[wall_11,floor_203]=True
    close[wall_11,wall_211]=True
    close[wall_11,ceiling_216]=True
    close[wall_11,cupboard_229]=True
    close[wall_11,kitchen_counter_230]=True
    close[wall_11,sink_231]=True
    close[wall_11,faucet_232]=True
    close[wall_11,fridge_289]=True
    close[wall_11,coffe_maker_290]=True
    close[wall_11,toaster_292]=True
    close[wall_11,microwave_297]=True
    close[wall_12,floor_2]=True
    close[wall_12,floor_3]=True
    close[wall_12,floor_4]=True
    close[wall_12,floor_6]=True
    close[wall_12,wall_9]=True
    close[wall_12,wall_14]=True
    close[wall_12,ceiling_16]=True
    close[wall_12,ceiling_17]=True
    close[wall_12,ceiling_21]=True
    close[wall_12,mat_22]=True
    close[wall_12,ceilinglamp_26]=True
    close[wall_12,walllamp_28]=True
    close[wall_12,towel_rack_31]=True
    close[wall_12,towel_rack_32]=True
    close[wall_12,bathroom_cabinet_40]=True
    close[wall_12,bathroom_counter_41]=True
    close[wall_12,sink_42]=True
    close[wall_12,faucet_43]=True
    close[wall_12,door_44]=True
    close[wall_12,doorjamb_45]=True
    close[wall_12,light_64]=True
    close[wall_12,floor_72]=True
    close[wall_12,wall_79]=True
    close[wall_12,ceiling_90]=True
    close[wall_12,bookshelf_101]=True
    close[wall_12,drawing_176]=True
    close[wall_12,photoframe_185]=True
    close[wall_13,floor_5]=True
    close[wall_13,wall_9]=True
    close[wall_13,wall_10]=True
    close[wall_13,ceiling_20]=True
    close[wall_13,curtain_23]=True
    close[wall_13,curtain_24]=True
    close[wall_13,curtain_25]=True
    close[wall_13,bathtub_30]=True
    close[wall_13,towel_rack_33]=True
    close[wall_13,towel_rack_34]=True
    close[wall_13,wallshelf_35]=True
    close[wall_13,window_63]=True
    close[wall_14,floor_6]=True
    close[wall_14,wall_11]=True
    close[wall_14,wall_12]=True
    close[wall_14,ceiling_17]=True
    close[wall_14,mat_22]=True
    close[wall_14,towel_rack_31]=True
    close[wall_14,towel_rack_32]=True
    close[wall_14,door_44]=True
    close[wall_14,doorjamb_45]=True
    close[wall_14,light_64]=True
    close[wall_14,floor_77]=True
    close[wall_14,wall_79]=True
    close[wall_14,wall_85]=True
    close[wall_14,ceiling_95]=True
    close[wall_14,bookshelf_101]=True
    close[wall_14,drawing_174]=True
    close[wall_14,photoframe_185]=True
    close[wall_14,wall_211]=True
    close[wall_14,fridge_289]=True
    close[wall_14,microwave_297]=True
    close[wall_15,floor_7]=True
    close[wall_15,wall_11]=True
    close[wall_15,ceiling_18]=True
    close[wall_15,walllamp_29]=True
    close[wall_15,shower_36]=True
    close[wall_15,toilet_37]=True
    close[wall_15,curtain_39]=True
    close[wall_15,floor_204]=True
    close[wall_15,wall_212]=True
    close[wall_15,ceiling_221]=True
    close[wall_15,cupboard_229]=True
    close[wall_15,kitchen_counter_230]=True
    close[wall_15,sink_231]=True
    close[wall_15,faucet_232]=True
    close[wall_15,stovefan_288]=True
    close[wall_15,coffe_maker_290]=True
    close[wall_15,toaster_292]=True
    close[wall_15,oven_295]=True
    close[wall_15,tray_296]=True
    close[wall_15,microwave_297]=True
    close[ceiling_16,wall_9]=True
    close[ceiling_16,wall_12]=True
    close[ceiling_16,ceiling_17]=True
    close[ceiling_16,ceiling_21]=True
    close[ceiling_16,ceilinglamp_26]=True
    close[ceiling_16,walllamp_28]=True
    close[ceiling_16,towel_rack_31]=True
    close[ceiling_16,towel_rack_32]=True
    close[ceiling_16,bathroom_cabinet_40]=True
    close[ceiling_16,faucet_43]=True
    close[ceiling_16,light_64]=True
    close[ceiling_16,wall_79]=True
    close[ceiling_16,ceiling_90]=True
    close[ceiling_16,bookshelf_101]=True
    close[ceiling_16,drawing_176]=True
    close[ceiling_16,photoframe_185]=True
    close[ceiling_17,wall_11]=True
    close[ceiling_17,wall_12]=True
    close[ceiling_17,wall_14]=True
    close[ceiling_17,ceiling_16]=True
    close[ceiling_17,ceiling_18]=True
    close[ceiling_17,ceiling_20]=True
    close[ceiling_17,ceilinglamp_26]=True
    close[ceiling_17,towel_rack_32]=True
    close[ceiling_17,doorjamb_45]=True
    close[ceiling_17,light_64]=True
    close[ceiling_17,wall_85]=True
    close[ceiling_17,ceiling_95]=True
    close[ceiling_18,wall_10]=True
    close[ceiling_18,wall_11]=True
    close[ceiling_18,wall_15]=True
    close[ceiling_18,ceiling_17]=True
    close[ceiling_18,ceiling_19]=True
    close[ceiling_18,ceilinglamp_26]=True
    close[ceiling_18,walllamp_29]=True
    close[ceiling_18,shower_36]=True
    close[ceiling_18,wall_211]=True
    close[ceiling_18,ceiling_216]=True
    close[ceiling_18,cupboard_229]=True
    close[ceiling_18,faucet_232]=True
    close[ceiling_18,fridge_289]=True
    close[ceiling_18,microwave_297]=True
    close[ceiling_19,wall_10]=True
    close[ceiling_19,wall_11]=True
    close[ceiling_19,ceiling_18]=True
    close[ceiling_19,ceiling_20]=True
    close[ceiling_19,curtain_25]=True
    close[ceiling_19,ceilinglamp_26]=True
    close[ceiling_19,walllamp_29]=True
    close[ceiling_19,shower_38]=True
    close[ceiling_19,curtain_39]=True
    close[ceiling_20,wall_9]=True
    close[ceiling_20,wall_10]=True
    close[ceiling_20,wall_13]=True
    close[ceiling_20,ceiling_17]=True
    close[ceiling_20,ceiling_19]=True
    close[ceiling_20,ceiling_21]=True
    close[ceiling_20,curtain_23]=True
    close[ceiling_20,curtain_24]=True
    close[ceiling_20,curtain_25]=True
    close[ceiling_20,ceilinglamp_26]=True
    close[ceiling_20,towel_rack_33]=True
    close[ceiling_20,wallshelf_35]=True
    close[ceiling_20,window_63]=True
    close[ceiling_21,wall_9]=True
    close[ceiling_21,wall_12]=True
    close[ceiling_21,ceiling_16]=True
    close[ceiling_21,ceiling_20]=True
    close[ceiling_21,curtain_23]=True
    close[ceiling_21,curtain_24]=True
    close[ceiling_21,ceilinglamp_26]=True
    close[ceiling_21,walllamp_27]=True
    close[ceiling_21,towel_rack_33]=True
    close[ceiling_21,towel_rack_34]=True
    close[ceiling_21,wallshelf_35]=True
    close[ceiling_21,bathroom_cabinet_40]=True
    close[ceiling_21,faucet_43]=True
    close[mat_22,basket_for_clothes_2006]=True
    close[mat_22,floor_2]=True
    close[mat_22,floor_3]=True
    close[mat_22,floor_5]=True
    close[mat_22,floor_6]=True
    close[mat_22,floor_7]=True
    close[mat_22,wall_11]=True
    close[mat_22,wall_12]=True
    close[mat_22,wall_14]=True
    close[mat_22,door_44]=True
    close[mat_22,doorjamb_45]=True
    close[mat_22,light_64]=True
    close[mat_22,floor_77]=True
    close[mat_22,wall_85]=True
    close[mat_22,fridge_289]=True
    close[curtain_23,floor_5]=True
    close[curtain_23,wall_9]=True
    close[curtain_23,wall_13]=True
    close[curtain_23,ceiling_20]=True
    close[curtain_23,ceiling_21]=True
    close[curtain_23,curtain_24]=True
    close[curtain_23,curtain_25]=True
    close[curtain_23,bathtub_30]=True
    close[curtain_23,towel_rack_33]=True
    close[curtain_23,wallshelf_35]=True
    close[curtain_23,window_63]=True
    close[curtain_24,floor_5]=True
    close[curtain_24,wall_9]=True
    close[curtain_24,wall_13]=True
    close[curtain_24,ceiling_20]=True
    close[curtain_24,ceiling_21]=True
    close[curtain_24,curtain_23]=True
    close[curtain_24,curtain_25]=True
    close[curtain_24,bathtub_30]=True
    close[curtain_24,towel_rack_33]=True
    close[curtain_24,wallshelf_35]=True
    close[curtain_24,window_63]=True
    close[curtain_25,floor_5]=True
    close[curtain_25,wall_10]=True
    close[curtain_25,wall_13]=True
    close[curtain_25,ceiling_19]=True
    close[curtain_25,ceiling_20]=True
    close[curtain_25,curtain_23]=True
    close[curtain_25,curtain_24]=True
    close[curtain_25,bathtub_30]=True
    close[curtain_25,window_63]=True
    close[ceilinglamp_26,wall_9]=True
    close[ceilinglamp_26,wall_10]=True
    close[ceilinglamp_26,wall_11]=True
    close[ceilinglamp_26,wall_12]=True
    close[ceilinglamp_26,ceiling_16]=True
    close[ceilinglamp_26,ceiling_17]=True
    close[ceilinglamp_26,ceiling_18]=True
    close[ceilinglamp_26,ceiling_19]=True
    close[ceilinglamp_26,ceiling_20]=True
    close[ceilinglamp_26,ceiling_21]=True
    close[walllamp_27,floor_4]=True
    close[walllamp_27,wall_9]=True
    close[walllamp_27,ceiling_21]=True
    close[walllamp_27,towel_rack_34]=True
    close[walllamp_27,wallshelf_35]=True
    close[walllamp_27,bathroom_cabinet_40]=True
    close[walllamp_27,bathroom_counter_41]=True
    close[walllamp_28,floor_2]=True
    close[walllamp_28,floor_3]=True
    close[walllamp_28,wall_12]=True
    close[walllamp_28,ceiling_16]=True
    close[walllamp_28,towel_rack_31]=True
    close[walllamp_28,towel_rack_32]=True
    close[walllamp_28,bathroom_cabinet_40]=True
    close[walllamp_28,bathroom_counter_41]=True
    close[walllamp_28,floor_71]=True
    close[walllamp_28,floor_72]=True
    close[walllamp_28,wall_79]=True
    close[walllamp_28,wall_82]=True
    close[walllamp_28,ceiling_89]=True
    close[walllamp_28,ceiling_90]=True
    close[walllamp_28,bookshelf_101]=True
    close[walllamp_28,drawing_176]=True
    close[walllamp_28,photoframe_185]=True
    close[walllamp_29,floor_7]=True
    close[walllamp_29,floor_8]=True
    close[walllamp_29,wall_10]=True
    close[walllamp_29,wall_11]=True
    close[walllamp_29,wall_15]=True
    close[walllamp_29,ceiling_18]=True
    close[walllamp_29,ceiling_19]=True
    close[walllamp_29,shower_36]=True
    close[walllamp_29,shower_38]=True
    close[walllamp_29,curtain_39]=True
    close[bathtub_30,basket_for_clothes_2006]=True
    close[bathtub_30,floor_4]=True
    close[bathtub_30,floor_5]=True
    close[bathtub_30,floor_8]=True
    close[bathtub_30,wall_9]=True
    close[bathtub_30,wall_10]=True
    close[bathtub_30,wall_13]=True
    close[bathtub_30,curtain_23]=True
    close[bathtub_30,curtain_24]=True
    close[bathtub_30,curtain_25]=True
    close[bathtub_30,towel_rack_33]=True
    close[bathtub_30,wallshelf_35]=True
    close[bathtub_30,window_63]=True
    close[towel_rack_31,basket_for_clothes_2006]=True
    close[towel_rack_31,towel_2056]=True
    close[towel_rack_31,floor_2]=True
    close[towel_rack_31,floor_3]=True
    close[towel_rack_31,wall_12]=True
    close[towel_rack_31,wall_14]=True
    close[towel_rack_31,ceiling_16]=True
    close[towel_rack_31,walllamp_28]=True
    close[towel_rack_31,towel_rack_32]=True
    close[towel_rack_31,bathroom_cabinet_40]=True
    close[towel_rack_31,bathroom_counter_41]=True
    close[towel_rack_31,floor_72]=True
    close[towel_rack_31,wall_79]=True
    close[towel_rack_31,wall_82]=True
    close[towel_rack_31,wall_85]=True
    close[towel_rack_31,ceiling_90]=True
    close[towel_rack_31,bookshelf_101]=True
    close[towel_rack_31,drawing_176]=True
    close[towel_rack_31,photoframe_185]=True
    close[towel_rack_32,basket_for_clothes_2006]=True
    close[towel_rack_32,towel_2057]=True
    close[towel_rack_32,floor_2]=True
    close[towel_rack_32,floor_3]=True
    close[towel_rack_32,floor_6]=True
    close[towel_rack_32,wall_12]=True
    close[towel_rack_32,wall_14]=True
    close[towel_rack_32,ceiling_16]=True
    close[towel_rack_32,ceiling_17]=True
    close[towel_rack_32,walllamp_28]=True
    close[towel_rack_32,towel_rack_31]=True
    close[towel_rack_32,bathroom_counter_41]=True
    close[towel_rack_32,light_64]=True
    close[towel_rack_32,floor_72]=True
    close[towel_rack_32,floor_77]=True
    close[towel_rack_32,wall_79]=True
    close[towel_rack_32,wall_85]=True
    close[towel_rack_32,ceiling_90]=True
    close[towel_rack_32,ceiling_95]=True
    close[towel_rack_32,bookshelf_101]=True
    close[towel_rack_32,photoframe_185]=True
    close[towel_rack_33,basket_for_clothes_2006]=True
    close[towel_rack_33,towel_2058]=True
    close[towel_rack_33,floor_4]=True
    close[towel_rack_33,floor_5]=True
    close[towel_rack_33,wall_9]=True
    close[towel_rack_33,wall_13]=True
    close[towel_rack_33,ceiling_20]=True
    close[towel_rack_33,ceiling_21]=True
    close[towel_rack_33,curtain_23]=True
    close[towel_rack_33,curtain_24]=True
    close[towel_rack_33,bathtub_30]=True
    close[towel_rack_33,towel_rack_34]=True
    close[towel_rack_33,wallshelf_35]=True
    close[towel_rack_33,window_63]=True
    close[towel_rack_34,basket_for_clothes_2006]=True
    close[towel_rack_34,towel_2059]=True
    close[towel_rack_34,floor_4]=True
    close[towel_rack_34,wall_9]=True
    close[towel_rack_34,wall_13]=True
    close[towel_rack_34,ceiling_21]=True
    close[towel_rack_34,walllamp_27]=True
    close[towel_rack_34,towel_rack_33]=True
    close[towel_rack_34,wallshelf_35]=True
    close[towel_rack_34,bathroom_counter_41]=True
    close[wallshelf_35,wall_9]=True
    close[wallshelf_35,wall_13]=True
    close[wallshelf_35,ceiling_20]=True
    close[wallshelf_35,ceiling_21]=True
    close[wallshelf_35,curtain_23]=True
    close[wallshelf_35,curtain_24]=True
    close[wallshelf_35,walllamp_27]=True
    close[wallshelf_35,bathtub_30]=True
    close[wallshelf_35,towel_rack_33]=True
    close[wallshelf_35,towel_rack_34]=True
    close[shower_36,basket_for_clothes_2006]=True
    close[shower_36,floor_7]=True
    close[shower_36,wall_11]=True
    close[shower_36,wall_15]=True
    close[shower_36,ceiling_18]=True
    close[shower_36,walllamp_29]=True
    close[shower_36,toilet_37]=True
    close[shower_36,floor_202]=True
    close[shower_36,floor_203]=True
    close[shower_36,wall_211]=True
    close[shower_36,wall_212]=True
    close[shower_36,ceiling_216]=True
    close[shower_36,cupboard_229]=True
    close[shower_36,kitchen_counter_230]=True
    close[shower_36,sink_231]=True
    close[shower_36,faucet_232]=True
    close[shower_36,fridge_289]=True
    close[shower_36,coffe_maker_290]=True
    close[shower_36,toaster_292]=True
    close[shower_36,microwave_297]=True
    close[toilet_37,basket_for_clothes_2006]=True
    close[toilet_37,floor_7]=True
    close[toilet_37,wall_11]=True
    close[toilet_37,wall_15]=True
    close[toilet_37,shower_36]=True
    close[toilet_37,floor_202]=True
    close[toilet_37,floor_203]=True
    close[toilet_37,floor_204]=True
    close[toilet_37,wall_211]=True
    close[toilet_37,wall_212]=True
    close[toilet_37,kitchen_counter_230]=True
    close[toilet_37,sink_231]=True
    close[toilet_37,faucet_232]=True
    close[toilet_37,fridge_289]=True
    close[toilet_37,toaster_292]=True
    close[toilet_37,microwave_297]=True
    close[shower_38,floor_8]=True
    close[shower_38,wall_10]=True
    close[shower_38,ceiling_19]=True
    close[shower_38,walllamp_29]=True
    close[shower_38,curtain_39]=True
    close[curtain_39,floor_8]=True
    close[curtain_39,wall_10]=True
    close[curtain_39,wall_11]=True
    close[curtain_39,wall_15]=True
    close[curtain_39,ceiling_19]=True
    close[curtain_39,walllamp_29]=True
    close[curtain_39,shower_38]=True
    close[bathroom_cabinet_40,wall_9]=True
    close[bathroom_cabinet_40,wall_12]=True
    close[bathroom_cabinet_40,ceiling_16]=True
    close[bathroom_cabinet_40,ceiling_21]=True
    close[bathroom_cabinet_40,walllamp_27]=True
    close[bathroom_cabinet_40,walllamp_28]=True
    close[bathroom_cabinet_40,towel_rack_31]=True
    close[bathroom_cabinet_40,bathroom_counter_41]=True
    close[bathroom_cabinet_40,sink_42]=True
    close[bathroom_cabinet_40,faucet_43]=True
    close[bathroom_cabinet_40,drawing_176]=True
    close[bathroom_counter_41,floor_2]=True
    close[bathroom_counter_41,floor_3]=True
    close[bathroom_counter_41,floor_4]=True
    close[bathroom_counter_41,wall_9]=True
    close[bathroom_counter_41,wall_12]=True
    close[bathroom_counter_41,walllamp_27]=True
    close[bathroom_counter_41,walllamp_28]=True
    close[bathroom_counter_41,towel_rack_31]=True
    close[bathroom_counter_41,towel_rack_32]=True
    close[bathroom_counter_41,towel_rack_34]=True
    close[bathroom_counter_41,bathroom_cabinet_40]=True
    close[bathroom_counter_41,sink_42]=True
    close[bathroom_counter_41,faucet_43]=True
    close[bathroom_counter_41,wall_79]=True
    close[bathroom_counter_41,bookshelf_101]=True
    close[bathroom_counter_41,drawing_176]=True
    close[sink_42,basket_for_clothes_2006]=True
    close[sink_42,washing_machine_2007]=True
    close[sink_42,soap_2053]=True
    close[sink_42,cleaning_solution_2073]=True
    close[sink_42,detergent_2084]=True
    close[sink_42,floor_2]=True
    close[sink_42,floor_3]=True
    close[sink_42,floor_4]=True
    close[sink_42,wall_9]=True
    close[sink_42,wall_12]=True
    close[sink_42,bathroom_cabinet_40]=True
    close[sink_42,bathroom_counter_41]=True
    close[sink_42,faucet_43]=True
    close[faucet_43,basket_for_clothes_2006]=True
    close[faucet_43,floor_2]=True
    close[faucet_43,floor_3]=True
    close[faucet_43,floor_4]=True
    close[faucet_43,wall_9]=True
    close[faucet_43,wall_12]=True
    close[faucet_43,ceiling_16]=True
    close[faucet_43,ceiling_21]=True
    close[faucet_43,bathroom_cabinet_40]=True
    close[faucet_43,bathroom_counter_41]=True
    close[faucet_43,sink_42]=True
    close[door_44,floor_2]=True
    close[door_44,floor_3]=True
    close[door_44,floor_6]=True
    close[door_44,floor_7]=True
    close[door_44,wall_11]=True
    close[door_44,wall_12]=True
    close[door_44,wall_14]=True
    close[door_44,mat_22]=True
    close[door_44,doorjamb_45]=True
    close[door_44,light_64]=True
    close[door_44,floor_72]=True
    close[door_44,floor_77]=True
    close[door_44,wall_79]=True
    close[door_44,wall_85]=True
    close[door_44,bookshelf_101]=True
    close[door_44,drawing_174]=True
    close[door_44,floor_202]=True
    close[door_44,floor_203]=True
    close[door_44,wall_211]=True
    close[door_44,fridge_289]=True
    close[doorjamb_45,floor_6]=True
    close[doorjamb_45,wall_11]=True
    close[doorjamb_45,wall_12]=True
    close[doorjamb_45,wall_14]=True
    close[doorjamb_45,ceiling_17]=True
    close[doorjamb_45,mat_22]=True
    close[doorjamb_45,door_44]=True
    close[doorjamb_45,light_64]=True
    close[doorjamb_45,floor_77]=True
    close[doorjamb_45,wall_79]=True
    close[doorjamb_45,wall_85]=True
    close[doorjamb_45,ceiling_95]=True
    close[doorjamb_45,bookshelf_101]=True
    close[doorjamb_45,drawing_174]=True
    close[doorjamb_45,wall_211]=True
    close[doorjamb_45,fridge_289]=True
    close[window_63,floor_5]=True
    close[window_63,wall_9]=True
    close[window_63,wall_10]=True
    close[window_63,wall_13]=True
    close[window_63,ceiling_20]=True
    close[window_63,curtain_23]=True
    close[window_63,curtain_24]=True
    close[window_63,curtain_25]=True
    close[window_63,bathtub_30]=True
    close[window_63,towel_rack_33]=True
    close[light_64,floor_2]=True
    close[light_64,floor_3]=True
    close[light_64,floor_6]=True
    close[light_64,wall_12]=True
    close[light_64,wall_14]=True
    close[light_64,ceiling_16]=True
    close[light_64,ceiling_17]=True
    close[light_64,mat_22]=True
    close[light_64,towel_rack_32]=True
    close[light_64,door_44]=True
    close[light_64,doorjamb_45]=True
    close[light_64,floor_72]=True
    close[light_64,floor_77]=True
    close[light_64,wall_79]=True
    close[light_64,wall_85]=True
    close[light_64,ceiling_90]=True
    close[light_64,ceiling_95]=True
    close[light_64,bookshelf_101]=True
    close[floor_68,floor_69]=True
    close[floor_68,floor_70]=True
    close[floor_68,floor_74]=True
    close[floor_68,wall_81]=True
    close[floor_68,tablelamp_97]=True
    close[floor_68,nightstand_100]=True
    close[floor_68,bed_105]=True
    close[floor_68,dresser_108]=True
    close[floor_68,closetdrawer_116]=True
    close[floor_68,closetdrawer_117]=True
    close[floor_68,closetdrawer_118]=True
    close[floor_68,closetdrawer_119]=True
    close[floor_68,closetdrawer_120]=True
    close[floor_68,closetdrawer_121]=True
    close[floor_68,closetdrawer_122]=True
    close[floor_68,dresser_123]=True
    close[floor_68,closetdrawer_143]=True
    close[floor_68,closetdrawer_146]=True
    close[floor_68,closetdrawer_148]=True
    close[floor_68,closetdrawer_150]=True
    close[floor_68,closetdrawer_154]=True
    close[floor_68,closetdrawer_158]=True
    close[floor_68,closetdrawer_160]=True
    close[floor_68,mat_173]=True
    close[floor_68,pillow_183]=True
    close[floor_69,floor_68]=True
    close[floor_69,floor_70]=True
    close[floor_69,floor_74]=True
    close[floor_69,wall_81]=True
    close[floor_69,tablelamp_97]=True
    close[floor_69,nightstand_100]=True
    close[floor_69,bed_105]=True
    close[floor_69,dresser_108]=True
    close[floor_69,closetdrawer_116]=True
    close[floor_69,closetdrawer_117]=True
    close[floor_69,closetdrawer_118]=True
    close[floor_69,closetdrawer_119]=True
    close[floor_69,closetdrawer_120]=True
    close[floor_69,closetdrawer_121]=True
    close[floor_69,closetdrawer_122]=True
    close[floor_69,dresser_123]=True
    close[floor_69,closetdrawer_143]=True
    close[floor_69,closetdrawer_146]=True
    close[floor_69,closetdrawer_148]=True
    close[floor_69,closetdrawer_150]=True
    close[floor_69,closetdrawer_154]=True
    close[floor_69,closetdrawer_158]=True
    close[floor_69,closetdrawer_160]=True
    close[floor_69,mat_173]=True
    close[floor_69,pillow_183]=True
    close[floor_69,chair_2004]=True
    close[floor_70,floor_68]=True
    close[floor_70,floor_69]=True
    close[floor_70,floor_71]=True
    close[floor_70,floor_73]=True
    close[floor_70,wall_80]=True
    close[floor_70,wall_81]=True
    close[floor_70,wall_82]=True
    close[floor_70,window_86]=True
    close[floor_70,tablelamp_97]=True
    close[floor_70,tablelamp_98]=True
    close[floor_70,nightstand_100]=True
    close[floor_70,nightstand_102]=True
    close[floor_70,bed_105]=True
    close[floor_70,mat_173]=True
    close[floor_70,curtain_179]=True
    close[floor_70,curtain_180]=True
    close[floor_70,curtain_181]=True
    close[floor_70,pillow_182]=True
    close[floor_70,pillow_183]=True
    close[floor_71,walllamp_28]=True
    close[floor_71,floor_70]=True
    close[floor_71,floor_72]=True
    close[floor_71,wall_82]=True
    close[floor_71,tablelamp_98]=True
    close[floor_71,nightstand_102]=True
    close[floor_71,bed_105]=True
    close[floor_71,chair_106]=True
    close[floor_71,mat_173]=True
    close[floor_71,drawing_176]=True
    close[floor_71,pillow_182]=True
    close[floor_72,floor_2]=True
    close[floor_72,floor_3]=True
    close[floor_72,wall_12]=True
    close[floor_72,walllamp_28]=True
    close[floor_72,towel_rack_31]=True
    close[floor_72,towel_rack_32]=True
    close[floor_72,door_44]=True
    close[floor_72,light_64]=True
    close[floor_72,floor_71]=True
    close[floor_72,floor_73]=True
    close[floor_72,floor_77]=True
    close[floor_72,wall_79]=True
    close[floor_72,wall_82]=True
    close[floor_72,wall_85]=True
    close[floor_72,bookshelf_101]=True
    close[floor_72,table_107]=True
    close[floor_72,mat_173]=True
    close[floor_72,orchid_178]=True
    close[floor_73,floor_70]=True
    close[floor_73,floor_72]=True
    close[floor_73,floor_74]=True
    close[floor_73,floor_76]=True
    close[floor_73,bed_105]=True
    close[floor_73,table_107]=True
    close[floor_73,mat_173]=True
    close[floor_73,orchid_178]=True
    close[floor_74,floor_68]=True
    close[floor_74,floor_69]=True
    close[floor_74,floor_73]=True
    close[floor_74,floor_75]=True
    close[floor_74,wall_78]=True
    close[floor_74,wall_81]=True
    close[floor_74,wall_83]=True
    close[floor_74,table_107]=True
    close[floor_74,dresser_108]=True
    close[floor_74,closetdrawer_116]=True
    close[floor_74,closetdrawer_117]=True
    close[floor_74,closetdrawer_118]=True
    close[floor_74,closetdrawer_119]=True
    close[floor_74,closetdrawer_120]=True
    close[floor_74,closetdrawer_121]=True
    close[floor_74,closetdrawer_122]=True
    close[floor_74,closetdrawer_154]=True
    close[floor_74,closetdrawer_160]=True
    close[floor_74,mat_173]=True
    close[floor_74,drawing_175]=True
    close[floor_74,orchid_178]=True
    close[floor_75,floor_74]=True
    close[floor_75,floor_76]=True
    close[floor_75,wall_83]=True
    close[floor_75,chair_103]=True
    close[floor_75,desk_104]=True
    close[floor_75,mouse_166]=True
    close[floor_75,mousepad_167]=True
    close[floor_75,keyboard_168]=True
    close[floor_75,light_169]=True
    close[floor_75,computer_170]=True
    close[floor_75,cpuscreen_171]=True
    close[floor_75,drawing_175]=True
    close[floor_75,floor_207]=True
    close[floor_75,wall_210]=True
    close[floor_75,door_222]=True
    close[floor_75,bookshelf_233]=True
    close[floor_76,floor_73]=True
    close[floor_76,floor_75]=True
    close[floor_76,floor_77]=True
    close[floor_76,wall_83]=True
    close[floor_76,wall_84]=True
    close[floor_76,wall_85]=True
    close[floor_76,trashcan_99]=True
    close[floor_76,chair_103]=True
    close[floor_76,desk_104]=True
    close[floor_76,table_107]=True
    close[floor_76,doorjamb_165]=True
    close[floor_76,keyboard_168]=True
    close[floor_76,light_169]=True
    close[floor_76,computer_170]=True
    close[floor_76,cpuscreen_171]=True
    close[floor_76,drawing_174]=True
    close[floor_76,orchid_178]=True
    close[floor_76,floor_206]=True
    close[floor_76,wall_209]=True
    close[floor_76,door_222]=True
    close[floor_76,bookshelf_233]=True
    close[floor_76,drawing_238]=True
    close[floor_76,light_245]=True
    close[floor_76,powersocket_246]=True
    close[floor_76,phone_247]=True
    close[floor_77,floor_6]=True
    close[floor_77,wall_14]=True
    close[floor_77,mat_22]=True
    close[floor_77,towel_rack_32]=True
    close[floor_77,door_44]=True
    close[floor_77,doorjamb_45]=True
    close[floor_77,light_64]=True
    close[floor_77,floor_72]=True
    close[floor_77,floor_76]=True
    close[floor_77,wall_85]=True
    close[floor_77,trashcan_99]=True
    close[floor_77,drawing_174]=True
    close[floor_77,floor_202]=True
    close[floor_77,floor_203]=True
    close[floor_77,wall_211]=True
    close[floor_77,door_222]=True
    close[floor_77,drawing_238]=True
    close[floor_77,light_245]=True
    close[floor_77,powersocket_246]=True
    close[floor_77,phone_247]=True
    close[floor_77,fridge_289]=True
    close[wall_78,floor_74]=True
    close[wall_78,wall_81]=True
    close[wall_78,wall_83]=True
    close[wall_78,ceiling_92]=True
    close[wall_78,dresser_108]=True
    close[wall_78,hanger_109]=True
    close[wall_78,hanger_110]=True
    close[wall_78,hanger_111]=True
    close[wall_78,hanger_112]=True
    close[wall_78,hanger_113]=True
    close[wall_78,hanger_114]=True
    close[wall_78,hanger_115]=True
    close[wall_78,closetdrawer_116]=True
    close[wall_78,closetdrawer_117]=True
    close[wall_78,closetdrawer_118]=True
    close[wall_78,closetdrawer_119]=True
    close[wall_78,closetdrawer_120]=True
    close[wall_78,closetdrawer_121]=True
    close[wall_78,closetdrawer_122]=True
    close[wall_78,hanger_126]=True
    close[wall_78,hanger_130]=True
    close[wall_78,hanger_132]=True
    close[wall_78,hanger_134]=True
    close[wall_78,hanger_136]=True
    close[wall_78,closetdrawer_143]=True
    close[wall_78,closetdrawer_150]=True
    close[wall_78,closetdrawer_154]=True
    close[wall_78,closetdrawer_160]=True
    close[wall_78,drawing_175]=True
    close[wall_79,floor_2]=True
    close[wall_79,floor_3]=True
    close[wall_79,wall_12]=True
    close[wall_79,wall_14]=True
    close[wall_79,ceiling_16]=True
    close[wall_79,walllamp_28]=True
    close[wall_79,towel_rack_31]=True
    close[wall_79,towel_rack_32]=True
    close[wall_79,bathroom_counter_41]=True
    close[wall_79,door_44]=True
    close[wall_79,doorjamb_45]=True
    close[wall_79,light_64]=True
    close[wall_79,floor_72]=True
    close[wall_79,wall_82]=True
    close[wall_79,wall_85]=True
    close[wall_79,ceiling_90]=True
    close[wall_79,bookshelf_101]=True
    close[wall_79,drawing_176]=True
    close[wall_79,photoframe_185]=True
    close[wall_80,floor_70]=True
    close[wall_80,wall_81]=True
    close[wall_80,wall_82]=True
    close[wall_80,window_86]=True
    close[wall_80,ceiling_88]=True
    close[wall_80,tablelamp_97]=True
    close[wall_80,tablelamp_98]=True
    close[wall_80,nightstand_100]=True
    close[wall_80,nightstand_102]=True
    close[wall_80,bed_105]=True
    close[wall_80,mat_173]=True
    close[wall_80,curtain_179]=True
    close[wall_80,curtain_180]=True
    close[wall_80,curtain_181]=True
    close[wall_80,pillow_182]=True
    close[wall_80,pillow_183]=True
    close[wall_81,floor_68]=True
    close[wall_81,floor_69]=True
    close[wall_81,floor_70]=True
    close[wall_81,floor_74]=True
    close[wall_81,wall_78]=True
    close[wall_81,wall_80]=True
    close[wall_81,window_86]=True
    close[wall_81,ceiling_87]=True
    close[wall_81,ceiling_88]=True
    close[wall_81,ceiling_92]=True
    close[wall_81,tablelamp_97]=True
    close[wall_81,nightstand_100]=True
    close[wall_81,bed_105]=True
    close[wall_81,dresser_108]=True
    close[wall_81,hanger_109]=True
    close[wall_81,hanger_110]=True
    close[wall_81,hanger_111]=True
    close[wall_81,hanger_112]=True
    close[wall_81,hanger_113]=True
    close[wall_81,hanger_114]=True
    close[wall_81,hanger_115]=True
    close[wall_81,closetdrawer_116]=True
    close[wall_81,closetdrawer_117]=True
    close[wall_81,closetdrawer_118]=True
    close[wall_81,closetdrawer_119]=True
    close[wall_81,closetdrawer_120]=True
    close[wall_81,closetdrawer_121]=True
    close[wall_81,closetdrawer_122]=True
    close[wall_81,dresser_123]=True
    close[wall_81,hanger_124]=True
    close[wall_81,hanger_126]=True
    close[wall_81,hanger_128]=True
    close[wall_81,hanger_130]=True
    close[wall_81,hanger_132]=True
    close[wall_81,hanger_134]=True
    close[wall_81,hanger_136]=True
    close[wall_81,hanger_138]=True
    close[wall_81,hanger_140]=True
    close[wall_81,hanger_141]=True
    close[wall_81,hanger_142]=True
    close[wall_81,closetdrawer_143]=True
    close[wall_81,closetdrawer_146]=True
    close[wall_81,closetdrawer_148]=True
    close[wall_81,closetdrawer_150]=True
    close[wall_81,closetdrawer_154]=True
    close[wall_81,closetdrawer_158]=True
    close[wall_81,closetdrawer_160]=True
    close[wall_81,mat_173]=True
    close[wall_81,curtain_179]=True
    close[wall_81,curtain_180]=True
    close[wall_81,pillow_183]=True
    close[wall_82,walllamp_28]=True
    close[wall_82,towel_rack_31]=True
    close[wall_82,floor_70]=True
    close[wall_82,floor_71]=True
    close[wall_82,floor_72]=True
    close[wall_82,wall_79]=True
    close[wall_82,wall_80]=True
    close[wall_82,window_86]=True
    close[wall_82,ceiling_88]=True
    close[wall_82,ceiling_89]=True
    close[wall_82,ceiling_90]=True
    close[wall_82,tablelamp_98]=True
    close[wall_82,bookshelf_101]=True
    close[wall_82,nightstand_102]=True
    close[wall_82,bed_105]=True
    close[wall_82,chair_106]=True
    close[wall_82,mat_173]=True
    close[wall_82,drawing_176]=True
    close[wall_82,curtain_181]=True
    close[wall_82,pillow_182]=True
    close[wall_82,photoframe_185]=True
    close[wall_83,floor_74]=True
    close[wall_83,floor_75]=True
    close[wall_83,floor_76]=True
    close[wall_83,wall_78]=True
    close[wall_83,wall_84]=True
    close[wall_83,ceiling_92]=True
    close[wall_83,ceiling_93]=True
    close[wall_83,ceiling_94]=True
    close[wall_83,chair_103]=True
    close[wall_83,desk_104]=True
    close[wall_83,doorjamb_165]=True
    close[wall_83,mouse_166]=True
    close[wall_83,mousepad_167]=True
    close[wall_83,keyboard_168]=True
    close[wall_83,light_169]=True
    close[wall_83,computer_170]=True
    close[wall_83,cpuscreen_171]=True
    close[wall_83,drawing_175]=True
    close[wall_83,floor_207]=True
    close[wall_83,wall_209]=True
    close[wall_83,wall_210]=True
    close[wall_83,ceiling_218]=True
    close[wall_83,door_222]=True
    close[wall_83,bookshelf_233]=True
    close[wall_84,floor_76]=True
    close[wall_84,wall_83]=True
    close[wall_84,wall_85]=True
    close[wall_84,ceiling_94]=True
    close[wall_84,trashcan_99]=True
    close[wall_84,chair_103]=True
    close[wall_84,desk_104]=True
    close[wall_84,doorjamb_165]=True
    close[wall_84,keyboard_168]=True
    close[wall_84,light_169]=True
    close[wall_84,computer_170]=True
    close[wall_84,cpuscreen_171]=True
    close[wall_84,drawing_174]=True
    close[wall_84,floor_206]=True
    close[wall_84,wall_209]=True
    close[wall_84,wall_210]=True
    close[wall_84,wall_211]=True
    close[wall_84,ceiling_217]=True
    close[wall_84,door_222]=True
    close[wall_84,bookshelf_233]=True
    close[wall_84,drawing_238]=True
    close[wall_84,drawing_239]=True
    close[wall_84,drawing_240]=True
    close[wall_84,light_245]=True
    close[wall_84,powersocket_246]=True
    close[wall_84,phone_247]=True
    close[wall_84,wall_clock_249]=True
    close[wall_85,floor_6]=True
    close[wall_85,wall_14]=True
    close[wall_85,ceiling_17]=True
    close[wall_85,mat_22]=True
    close[wall_85,towel_rack_31]=True
    close[wall_85,towel_rack_32]=True
    close[wall_85,door_44]=True
    close[wall_85,doorjamb_45]=True
    close[wall_85,light_64]=True
    close[wall_85,floor_72]=True
    close[wall_85,floor_76]=True
    close[wall_85,floor_77]=True
    close[wall_85,wall_79]=True
    close[wall_85,wall_84]=True
    close[wall_85,ceiling_90]=True
    close[wall_85,ceiling_94]=True
    close[wall_85,ceiling_95]=True
    close[wall_85,trashcan_99]=True
    close[wall_85,bookshelf_101]=True
    close[wall_85,doorjamb_165]=True
    close[wall_85,drawing_174]=True
    close[wall_85,photoframe_185]=True
    close[wall_85,floor_202]=True
    close[wall_85,floor_203]=True
    close[wall_85,wall_209]=True
    close[wall_85,wall_211]=True
    close[wall_85,ceiling_216]=True
    close[wall_85,door_222]=True
    close[wall_85,drawing_238]=True
    close[wall_85,drawing_239]=True
    close[wall_85,drawing_240]=True
    close[wall_85,light_245]=True
    close[wall_85,powersocket_246]=True
    close[wall_85,phone_247]=True
    close[wall_85,wall_clock_249]=True
    close[wall_85,fridge_289]=True
    close[wall_85,microwave_297]=True
    close[window_86,floor_70]=True
    close[window_86,wall_80]=True
    close[window_86,wall_81]=True
    close[window_86,wall_82]=True
    close[window_86,ceiling_88]=True
    close[window_86,tablelamp_97]=True
    close[window_86,tablelamp_98]=True
    close[window_86,nightstand_100]=True
    close[window_86,nightstand_102]=True
    close[window_86,bed_105]=True
    close[window_86,mat_173]=True
    close[window_86,curtain_179]=True
    close[window_86,curtain_180]=True
    close[window_86,curtain_181]=True
    close[window_86,pillow_182]=True
    close[window_86,pillow_183]=True
    close[ceiling_87,wall_81]=True
    close[ceiling_87,ceiling_88]=True
    close[ceiling_87,ceiling_92]=True
    close[ceiling_87,dresser_108]=True
    close[ceiling_87,hanger_109]=True
    close[ceiling_87,hanger_110]=True
    close[ceiling_87,hanger_111]=True
    close[ceiling_87,hanger_112]=True
    close[ceiling_87,hanger_113]=True
    close[ceiling_87,hanger_114]=True
    close[ceiling_87,hanger_115]=True
    close[ceiling_87,dresser_123]=True
    close[ceiling_87,hanger_124]=True
    close[ceiling_87,hanger_126]=True
    close[ceiling_87,hanger_128]=True
    close[ceiling_87,hanger_130]=True
    close[ceiling_87,hanger_132]=True
    close[ceiling_87,hanger_134]=True
    close[ceiling_87,hanger_136]=True
    close[ceiling_87,hanger_138]=True
    close[ceiling_87,hanger_140]=True
    close[ceiling_87,hanger_141]=True
    close[ceiling_87,hanger_142]=True
    close[ceiling_87,curtain_179]=True
    close[ceiling_87,curtain_180]=True
    close[ceiling_88,wall_80]=True
    close[ceiling_88,wall_81]=True
    close[ceiling_88,wall_82]=True
    close[ceiling_88,window_86]=True
    close[ceiling_88,ceiling_87]=True
    close[ceiling_88,ceiling_89]=True
    close[ceiling_88,ceiling_91]=True
    close[ceiling_88,ceilinglamp_96]=True
    close[ceiling_88,curtain_179]=True
    close[ceiling_88,curtain_180]=True
    close[ceiling_88,curtain_181]=True
    close[ceiling_89,walllamp_28]=True
    close[ceiling_89,wall_82]=True
    close[ceiling_89,ceiling_88]=True
    close[ceiling_89,ceiling_90]=True
    close[ceiling_89,drawing_176]=True
    close[ceiling_89,curtain_181]=True
    close[ceiling_89,photoframe_185]=True
    close[ceiling_90,wall_12]=True
    close[ceiling_90,ceiling_16]=True
    close[ceiling_90,walllamp_28]=True
    close[ceiling_90,towel_rack_31]=True
    close[ceiling_90,towel_rack_32]=True
    close[ceiling_90,light_64]=True
    close[ceiling_90,wall_79]=True
    close[ceiling_90,wall_82]=True
    close[ceiling_90,wall_85]=True
    close[ceiling_90,ceiling_89]=True
    close[ceiling_90,ceiling_91]=True
    close[ceiling_90,ceiling_95]=True
    close[ceiling_90,ceilinglamp_96]=True
    close[ceiling_90,bookshelf_101]=True
    close[ceiling_90,photoframe_185]=True
    close[ceiling_91,ceiling_88]=True
    close[ceiling_91,ceiling_90]=True
    close[ceiling_91,ceiling_92]=True
    close[ceiling_91,ceiling_94]=True
    close[ceiling_91,ceilinglamp_96]=True
    close[ceiling_92,wall_78]=True
    close[ceiling_92,wall_81]=True
    close[ceiling_92,wall_83]=True
    close[ceiling_92,ceiling_87]=True
    close[ceiling_92,ceiling_91]=True
    close[ceiling_92,ceiling_93]=True
    close[ceiling_92,ceilinglamp_96]=True
    close[ceiling_92,dresser_108]=True
    close[ceiling_92,hanger_109]=True
    close[ceiling_92,hanger_110]=True
    close[ceiling_92,hanger_111]=True
    close[ceiling_92,hanger_112]=True
    close[ceiling_92,hanger_113]=True
    close[ceiling_92,hanger_114]=True
    close[ceiling_92,hanger_115]=True
    close[ceiling_92,hanger_126]=True
    close[ceiling_92,hanger_130]=True
    close[ceiling_92,hanger_132]=True
    close[ceiling_92,hanger_134]=True
    close[ceiling_92,drawing_175]=True
    close[ceiling_93,wall_83]=True
    close[ceiling_93,ceiling_92]=True
    close[ceiling_93,ceiling_94]=True
    close[ceiling_93,chair_103]=True
    close[ceiling_93,light_169]=True
    close[ceiling_93,cpuscreen_171]=True
    close[ceiling_93,drawing_175]=True
    close[ceiling_93,wall_210]=True
    close[ceiling_93,ceiling_218]=True
    close[ceiling_93,bookshelf_233]=True
    close[ceiling_94,wall_83]=True
    close[ceiling_94,wall_84]=True
    close[ceiling_94,wall_85]=True
    close[ceiling_94,ceiling_91]=True
    close[ceiling_94,ceiling_93]=True
    close[ceiling_94,ceiling_95]=True
    close[ceiling_94,ceilinglamp_96]=True
    close[ceiling_94,doorjamb_165]=True
    close[ceiling_94,light_169]=True
    close[ceiling_94,drawing_174]=True
    close[ceiling_94,wall_209]=True
    close[ceiling_94,ceiling_217]=True
    close[ceiling_94,drawing_238]=True
    close[ceiling_94,drawing_239]=True
    close[ceiling_94,drawing_240]=True
    close[ceiling_94,light_245]=True
    close[ceiling_94,phone_247]=True
    close[ceiling_94,wall_clock_249]=True
    close[ceiling_95,wall_14]=True
    close[ceiling_95,ceiling_17]=True
    close[ceiling_95,towel_rack_32]=True
    close[ceiling_95,doorjamb_45]=True
    close[ceiling_95,light_64]=True
    close[ceiling_95,wall_85]=True
    close[ceiling_95,ceiling_90]=True
    close[ceiling_95,ceiling_94]=True
    close[ceiling_95,drawing_174]=True
    close[ceiling_95,wall_211]=True
    close[ceiling_95,ceiling_216]=True
    close[ceiling_95,drawing_238]=True
    close[ceiling_95,drawing_239]=True
    close[ceiling_95,drawing_240]=True
    close[ceiling_95,light_245]=True
    close[ceiling_95,phone_247]=True
    close[ceiling_95,wall_clock_249]=True
    close[ceiling_95,fridge_289]=True
    close[ceilinglamp_96,ceiling_88]=True
    close[ceilinglamp_96,ceiling_90]=True
    close[ceilinglamp_96,ceiling_91]=True
    close[ceilinglamp_96,ceiling_92]=True
    close[ceilinglamp_96,ceiling_94]=True
    close[tablelamp_97,floor_68]=True
    close[tablelamp_97,floor_69]=True
    close[tablelamp_97,floor_70]=True
    close[tablelamp_97,wall_80]=True
    close[tablelamp_97,wall_81]=True
    close[tablelamp_97,window_86]=True
    close[tablelamp_97,nightstand_100]=True
    close[tablelamp_97,bed_105]=True
    close[tablelamp_97,mat_173]=True
    close[tablelamp_97,curtain_179]=True
    close[tablelamp_97,curtain_180]=True
    close[tablelamp_97,pillow_182]=True
    close[tablelamp_97,pillow_183]=True
    close[tablelamp_98,floor_70]=True
    close[tablelamp_98,floor_71]=True
    close[tablelamp_98,wall_80]=True
    close[tablelamp_98,wall_82]=True
    close[tablelamp_98,window_86]=True
    close[tablelamp_98,nightstand_102]=True
    close[tablelamp_98,bed_105]=True
    close[tablelamp_98,mat_173]=True
    close[tablelamp_98,curtain_181]=True
    close[tablelamp_98,pillow_182]=True
    close[tablelamp_98,pillow_183]=True
    close[trashcan_99,floor_76]=True
    close[trashcan_99,floor_77]=True
    close[trashcan_99,wall_84]=True
    close[trashcan_99,wall_85]=True
    close[trashcan_99,doorjamb_165]=True
    close[trashcan_99,drawing_174]=True
    close[trashcan_99,floor_202]=True
    close[trashcan_99,floor_203]=True
    close[trashcan_99,floor_206]=True
    close[trashcan_99,wall_209]=True
    close[trashcan_99,wall_211]=True
    close[trashcan_99,door_222]=True
    close[trashcan_99,kitchen_counter_230]=True
    close[trashcan_99,drawing_238]=True
    close[trashcan_99,drawing_239]=True
    close[trashcan_99,drawing_240]=True
    close[trashcan_99,light_245]=True
    close[trashcan_99,powersocket_246]=True
    close[trashcan_99,phone_247]=True
    close[trashcan_99,wall_clock_249]=True
    close[trashcan_99,fridge_289]=True
    close[nightstand_100,floor_68]=True
    close[nightstand_100,floor_69]=True
    close[nightstand_100,floor_70]=True
    close[nightstand_100,wall_80]=True
    close[nightstand_100,wall_81]=True
    close[nightstand_100,window_86]=True
    close[nightstand_100,tablelamp_97]=True
    close[nightstand_100,bed_105]=True
    close[nightstand_100,mat_173]=True
    close[nightstand_100,curtain_179]=True
    close[nightstand_100,curtain_180]=True
    close[nightstand_100,pillow_182]=True
    close[nightstand_100,pillow_183]=True
    close[bookshelf_101,floor_2]=True
    close[bookshelf_101,floor_3]=True
    close[bookshelf_101,wall_12]=True
    close[bookshelf_101,wall_14]=True
    close[bookshelf_101,ceiling_16]=True
    close[bookshelf_101,walllamp_28]=True
    close[bookshelf_101,towel_rack_31]=True
    close[bookshelf_101,towel_rack_32]=True
    close[bookshelf_101,bathroom_counter_41]=True
    close[bookshelf_101,door_44]=True
    close[bookshelf_101,doorjamb_45]=True
    close[bookshelf_101,light_64]=True
    close[bookshelf_101,floor_72]=True
    close[bookshelf_101,wall_79]=True
    close[bookshelf_101,wall_82]=True
    close[bookshelf_101,wall_85]=True
    close[bookshelf_101,ceiling_90]=True
    close[bookshelf_101,drawing_176]=True
    close[bookshelf_101,photoframe_185]=True
    close[nightstand_102,floor_70]=True
    close[nightstand_102,floor_71]=True
    close[nightstand_102,wall_80]=True
    close[nightstand_102,wall_82]=True
    close[nightstand_102,window_86]=True
    close[nightstand_102,tablelamp_98]=True
    close[nightstand_102,bed_105]=True
    close[nightstand_102,chair_106]=True
    close[nightstand_102,mat_173]=True
    close[nightstand_102,curtain_181]=True
    close[nightstand_102,pillow_182]=True
    close[nightstand_102,pillow_183]=True
    close[chair_103,floor_75]=True
    close[chair_103,floor_76]=True
    close[chair_103,wall_83]=True
    close[chair_103,wall_84]=True
    close[chair_103,ceiling_93]=True
    close[chair_103,desk_104]=True
    close[chair_103,mouse_166]=True
    close[chair_103,mousepad_167]=True
    close[chair_103,keyboard_168]=True
    close[chair_103,light_169]=True
    close[chair_103,computer_170]=True
    close[chair_103,cpuscreen_171]=True
    close[chair_103,floor_207]=True
    close[chair_103,wall_209]=True
    close[chair_103,wall_210]=True
    close[chair_103,bookshelf_233]=True
    close[desk_104,floor_75]=True
    close[desk_104,floor_76]=True
    close[desk_104,wall_83]=True
    close[desk_104,wall_84]=True
    close[desk_104,chair_103]=True
    close[desk_104,doorjamb_165]=True
    close[desk_104,mouse_166]=True
    close[desk_104,mousepad_167]=True
    close[desk_104,keyboard_168]=True
    close[desk_104,light_169]=True
    close[desk_104,computer_170]=True
    close[desk_104,cpuscreen_171]=True
    close[desk_104,drawing_175]=True
    close[desk_104,floor_206]=True
    close[desk_104,floor_207]=True
    close[desk_104,wall_209]=True
    close[desk_104,wall_210]=True
    close[desk_104,door_222]=True
    close[desk_104,bookshelf_233]=True
    close[bed_105,clothes_dress_2044]=True
    close[bed_105,clothes_scarf_2048]=True
    close[bed_105,clothes_underwear_2049]=True
    close[bed_105,floor_68]=True
    close[bed_105,floor_69]=True
    close[bed_105,floor_70]=True
    close[bed_105,floor_71]=True
    close[bed_105,floor_73]=True
    close[bed_105,wall_80]=True
    close[bed_105,wall_81]=True
    close[bed_105,wall_82]=True
    close[bed_105,window_86]=True
    close[bed_105,tablelamp_97]=True
    close[bed_105,tablelamp_98]=True
    close[bed_105,nightstand_100]=True
    close[bed_105,nightstand_102]=True
    close[bed_105,mat_173]=True
    close[bed_105,curtain_179]=True
    close[bed_105,curtain_180]=True
    close[bed_105,curtain_181]=True
    close[bed_105,pillow_182]=True
    close[bed_105,pillow_183]=True
    close[chair_106,floor_71]=True
    close[chair_106,wall_82]=True
    close[chair_106,nightstand_102]=True
    close[chair_106,mat_173]=True
    close[chair_106,drawing_176]=True
    close[table_107,clothes_hat_2045]=True
    close[table_107,clothes_gloves_2046]=True
    close[table_107,floor_72]=True
    close[table_107,floor_73]=True
    close[table_107,floor_74]=True
    close[table_107,floor_76]=True
    close[table_107,mat_173]=True
    close[table_107,orchid_178]=True
    close[dresser_108,floor_68]=True
    close[dresser_108,floor_69]=True
    close[dresser_108,floor_74]=True
    close[dresser_108,wall_78]=True
    close[dresser_108,wall_81]=True
    close[dresser_108,ceiling_87]=True
    close[dresser_108,ceiling_92]=True
    close[dresser_108,hanger_109]=True
    close[dresser_108,hanger_110]=True
    close[dresser_108,hanger_111]=True
    close[dresser_108,hanger_112]=True
    close[dresser_108,hanger_113]=True
    close[dresser_108,hanger_114]=True
    close[dresser_108,hanger_115]=True
    close[dresser_108,closetdrawer_116]=True
    close[dresser_108,closetdrawer_117]=True
    close[dresser_108,closetdrawer_118]=True
    close[dresser_108,closetdrawer_119]=True
    close[dresser_108,closetdrawer_120]=True
    close[dresser_108,closetdrawer_121]=True
    close[dresser_108,closetdrawer_122]=True
    close[dresser_108,dresser_123]=True
    close[dresser_108,hanger_124]=True
    close[dresser_108,hanger_126]=True
    close[dresser_108,hanger_128]=True
    close[dresser_108,hanger_130]=True
    close[dresser_108,hanger_132]=True
    close[dresser_108,hanger_134]=True
    close[dresser_108,hanger_136]=True
    close[dresser_108,hanger_138]=True
    close[dresser_108,hanger_140]=True
    close[dresser_108,hanger_141]=True
    close[dresser_108,hanger_142]=True
    close[dresser_108,closetdrawer_143]=True
    close[dresser_108,closetdrawer_146]=True
    close[dresser_108,closetdrawer_148]=True
    close[dresser_108,closetdrawer_150]=True
    close[dresser_108,closetdrawer_154]=True
    close[dresser_108,closetdrawer_158]=True
    close[dresser_108,closetdrawer_160]=True
    close[hanger_109,wall_78]=True
    close[hanger_109,wall_81]=True
    close[hanger_109,ceiling_87]=True
    close[hanger_109,ceiling_92]=True
    close[hanger_109,dresser_108]=True
    close[hanger_109,hanger_110]=True
    close[hanger_109,hanger_111]=True
    close[hanger_109,hanger_112]=True
    close[hanger_109,hanger_113]=True
    close[hanger_109,hanger_114]=True
    close[hanger_109,hanger_115]=True
    close[hanger_109,closetdrawer_116]=True
    close[hanger_109,closetdrawer_117]=True
    close[hanger_109,closetdrawer_118]=True
    close[hanger_109,closetdrawer_119]=True
    close[hanger_109,closetdrawer_120]=True
    close[hanger_109,dresser_123]=True
    close[hanger_109,hanger_126]=True
    close[hanger_109,hanger_128]=True
    close[hanger_109,hanger_130]=True
    close[hanger_109,hanger_132]=True
    close[hanger_109,hanger_134]=True
    close[hanger_109,hanger_136]=True
    close[hanger_109,hanger_138]=True
    close[hanger_109,closetdrawer_143]=True
    close[hanger_109,closetdrawer_150]=True
    close[hanger_109,closetdrawer_154]=True
    close[hanger_110,wall_78]=True
    close[hanger_110,wall_81]=True
    close[hanger_110,ceiling_87]=True
    close[hanger_110,ceiling_92]=True
    close[hanger_110,dresser_108]=True
    close[hanger_110,hanger_109]=True
    close[hanger_110,hanger_111]=True
    close[hanger_110,hanger_112]=True
    close[hanger_110,hanger_113]=True
    close[hanger_110,hanger_114]=True
    close[hanger_110,hanger_115]=True
    close[hanger_110,closetdrawer_116]=True
    close[hanger_110,closetdrawer_117]=True
    close[hanger_110,closetdrawer_118]=True
    close[hanger_110,closetdrawer_119]=True
    close[hanger_110,closetdrawer_120]=True
    close[hanger_110,dresser_123]=True
    close[hanger_110,hanger_126]=True
    close[hanger_110,hanger_128]=True
    close[hanger_110,hanger_130]=True
    close[hanger_110,hanger_132]=True
    close[hanger_110,hanger_134]=True
    close[hanger_110,hanger_136]=True
    close[hanger_110,hanger_138]=True
    close[hanger_110,closetdrawer_143]=True
    close[hanger_110,closetdrawer_150]=True
    close[hanger_111,wall_78]=True
    close[hanger_111,wall_81]=True
    close[hanger_111,ceiling_87]=True
    close[hanger_111,ceiling_92]=True
    close[hanger_111,dresser_108]=True
    close[hanger_111,hanger_109]=True
    close[hanger_111,hanger_110]=True
    close[hanger_111,hanger_112]=True
    close[hanger_111,hanger_113]=True
    close[hanger_111,hanger_114]=True
    close[hanger_111,hanger_115]=True
    close[hanger_111,closetdrawer_116]=True
    close[hanger_111,closetdrawer_117]=True
    close[hanger_111,closetdrawer_118]=True
    close[hanger_111,closetdrawer_119]=True
    close[hanger_111,closetdrawer_120]=True
    close[hanger_111,dresser_123]=True
    close[hanger_111,hanger_126]=True
    close[hanger_111,hanger_130]=True
    close[hanger_111,hanger_132]=True
    close[hanger_111,hanger_134]=True
    close[hanger_111,hanger_136]=True
    close[hanger_111,hanger_138]=True
    close[hanger_111,closetdrawer_143]=True
    close[hanger_111,closetdrawer_150]=True
    close[hanger_112,wall_78]=True
    close[hanger_112,wall_81]=True
    close[hanger_112,ceiling_87]=True
    close[hanger_112,ceiling_92]=True
    close[hanger_112,dresser_108]=True
    close[hanger_112,hanger_109]=True
    close[hanger_112,hanger_110]=True
    close[hanger_112,hanger_111]=True
    close[hanger_112,hanger_113]=True
    close[hanger_112,hanger_114]=True
    close[hanger_112,hanger_115]=True
    close[hanger_112,closetdrawer_116]=True
    close[hanger_112,closetdrawer_117]=True
    close[hanger_112,closetdrawer_118]=True
    close[hanger_112,closetdrawer_119]=True
    close[hanger_112,closetdrawer_120]=True
    close[hanger_112,dresser_123]=True
    close[hanger_112,hanger_126]=True
    close[hanger_112,hanger_130]=True
    close[hanger_112,hanger_132]=True
    close[hanger_112,hanger_134]=True
    close[hanger_112,hanger_136]=True
    close[hanger_112,closetdrawer_143]=True
    close[hanger_112,closetdrawer_150]=True
    close[hanger_113,wall_78]=True
    close[hanger_113,wall_81]=True
    close[hanger_113,ceiling_87]=True
    close[hanger_113,ceiling_92]=True
    close[hanger_113,dresser_108]=True
    close[hanger_113,hanger_109]=True
    close[hanger_113,hanger_110]=True
    close[hanger_113,hanger_111]=True
    close[hanger_113,hanger_112]=True
    close[hanger_113,hanger_114]=True
    close[hanger_113,hanger_115]=True
    close[hanger_113,closetdrawer_116]=True
    close[hanger_113,closetdrawer_117]=True
    close[hanger_113,closetdrawer_118]=True
    close[hanger_113,closetdrawer_119]=True
    close[hanger_113,closetdrawer_120]=True
    close[hanger_113,dresser_123]=True
    close[hanger_113,hanger_126]=True
    close[hanger_113,hanger_130]=True
    close[hanger_113,hanger_132]=True
    close[hanger_113,hanger_134]=True
    close[hanger_113,closetdrawer_143]=True
    close[hanger_114,wall_78]=True
    close[hanger_114,wall_81]=True
    close[hanger_114,ceiling_87]=True
    close[hanger_114,ceiling_92]=True
    close[hanger_114,dresser_108]=True
    close[hanger_114,hanger_109]=True
    close[hanger_114,hanger_110]=True
    close[hanger_114,hanger_111]=True
    close[hanger_114,hanger_112]=True
    close[hanger_114,hanger_113]=True
    close[hanger_114,hanger_115]=True
    close[hanger_114,closetdrawer_116]=True
    close[hanger_114,closetdrawer_117]=True
    close[hanger_114,closetdrawer_119]=True
    close[hanger_114,closetdrawer_120]=True
    close[hanger_114,dresser_123]=True
    close[hanger_114,hanger_132]=True
    close[hanger_115,wall_78]=True
    close[hanger_115,wall_81]=True
    close[hanger_115,ceiling_87]=True
    close[hanger_115,ceiling_92]=True
    close[hanger_115,dresser_108]=True
    close[hanger_115,hanger_109]=True
    close[hanger_115,hanger_110]=True
    close[hanger_115,hanger_111]=True
    close[hanger_115,hanger_112]=True
    close[hanger_115,hanger_113]=True
    close[hanger_115,hanger_114]=True
    close[hanger_115,closetdrawer_116]=True
    close[hanger_115,closetdrawer_117]=True
    close[hanger_115,closetdrawer_119]=True
    close[hanger_115,closetdrawer_120]=True
    close[hanger_115,dresser_123]=True
    close[hanger_115,hanger_126]=True
    close[hanger_115,hanger_132]=True
    close[hanger_115,hanger_134]=True
    close[closetdrawer_116,floor_68]=True
    close[closetdrawer_116,floor_69]=True
    close[closetdrawer_116,floor_74]=True
    close[closetdrawer_116,wall_78]=True
    close[closetdrawer_116,wall_81]=True
    close[closetdrawer_116,dresser_108]=True
    close[closetdrawer_116,hanger_109]=True
    close[closetdrawer_116,hanger_110]=True
    close[closetdrawer_116,hanger_111]=True
    close[closetdrawer_116,hanger_112]=True
    close[closetdrawer_116,hanger_113]=True
    close[closetdrawer_116,hanger_114]=True
    close[closetdrawer_116,hanger_115]=True
    close[closetdrawer_116,closetdrawer_117]=True
    close[closetdrawer_116,closetdrawer_118]=True
    close[closetdrawer_116,closetdrawer_119]=True
    close[closetdrawer_116,closetdrawer_120]=True
    close[closetdrawer_116,closetdrawer_121]=True
    close[closetdrawer_116,closetdrawer_122]=True
    close[closetdrawer_116,dresser_123]=True
    close[closetdrawer_116,hanger_126]=True
    close[closetdrawer_116,hanger_130]=True
    close[closetdrawer_116,hanger_132]=True
    close[closetdrawer_116,hanger_134]=True
    close[closetdrawer_116,hanger_136]=True
    close[closetdrawer_116,hanger_138]=True
    close[closetdrawer_116,closetdrawer_143]=True
    close[closetdrawer_116,closetdrawer_150]=True
    close[closetdrawer_116,closetdrawer_154]=True
    close[closetdrawer_116,closetdrawer_160]=True
    close[closetdrawer_117,floor_68]=True
    close[closetdrawer_117,floor_69]=True
    close[closetdrawer_117,floor_74]=True
    close[closetdrawer_117,wall_78]=True
    close[closetdrawer_117,wall_81]=True
    close[closetdrawer_117,dresser_108]=True
    close[closetdrawer_117,hanger_109]=True
    close[closetdrawer_117,hanger_110]=True
    close[closetdrawer_117,hanger_111]=True
    close[closetdrawer_117,hanger_112]=True
    close[closetdrawer_117,hanger_113]=True
    close[closetdrawer_117,hanger_114]=True
    close[closetdrawer_117,hanger_115]=True
    close[closetdrawer_117,closetdrawer_116]=True
    close[closetdrawer_117,closetdrawer_118]=True
    close[closetdrawer_117,closetdrawer_119]=True
    close[closetdrawer_117,closetdrawer_120]=True
    close[closetdrawer_117,closetdrawer_121]=True
    close[closetdrawer_117,closetdrawer_122]=True
    close[closetdrawer_117,dresser_123]=True
    close[closetdrawer_117,hanger_124]=True
    close[closetdrawer_117,hanger_126]=True
    close[closetdrawer_117,hanger_128]=True
    close[closetdrawer_117,hanger_130]=True
    close[closetdrawer_117,hanger_132]=True
    close[closetdrawer_117,hanger_134]=True
    close[closetdrawer_117,hanger_136]=True
    close[closetdrawer_117,hanger_138]=True
    close[closetdrawer_117,closetdrawer_143]=True
    close[closetdrawer_117,closetdrawer_146]=True
    close[closetdrawer_117,closetdrawer_148]=True
    close[closetdrawer_117,closetdrawer_150]=True
    close[closetdrawer_117,closetdrawer_154]=True
    close[closetdrawer_117,closetdrawer_158]=True
    close[closetdrawer_117,closetdrawer_160]=True
    close[closetdrawer_118,floor_68]=True
    close[closetdrawer_118,floor_69]=True
    close[closetdrawer_118,floor_74]=True
    close[closetdrawer_118,wall_78]=True
    close[closetdrawer_118,wall_81]=True
    close[closetdrawer_118,dresser_108]=True
    close[closetdrawer_118,hanger_109]=True
    close[closetdrawer_118,hanger_110]=True
    close[closetdrawer_118,hanger_111]=True
    close[closetdrawer_118,hanger_112]=True
    close[closetdrawer_118,hanger_113]=True
    close[closetdrawer_118,closetdrawer_116]=True
    close[closetdrawer_118,closetdrawer_117]=True
    close[closetdrawer_118,closetdrawer_119]=True
    close[closetdrawer_118,closetdrawer_120]=True
    close[closetdrawer_118,closetdrawer_121]=True
    close[closetdrawer_118,closetdrawer_122]=True
    close[closetdrawer_118,dresser_123]=True
    close[closetdrawer_118,hanger_126]=True
    close[closetdrawer_118,hanger_130]=True
    close[closetdrawer_118,hanger_132]=True
    close[closetdrawer_118,hanger_134]=True
    close[closetdrawer_118,hanger_136]=True
    close[closetdrawer_118,hanger_138]=True
    close[closetdrawer_118,closetdrawer_143]=True
    close[closetdrawer_118,closetdrawer_146]=True
    close[closetdrawer_118,closetdrawer_148]=True
    close[closetdrawer_118,closetdrawer_150]=True
    close[closetdrawer_118,closetdrawer_154]=True
    close[closetdrawer_118,closetdrawer_158]=True
    close[closetdrawer_118,closetdrawer_160]=True
    close[closetdrawer_119,floor_68]=True
    close[closetdrawer_119,floor_69]=True
    close[closetdrawer_119,floor_74]=True
    close[closetdrawer_119,wall_78]=True
    close[closetdrawer_119,wall_81]=True
    close[closetdrawer_119,dresser_108]=True
    close[closetdrawer_119,hanger_109]=True
    close[closetdrawer_119,hanger_110]=True
    close[closetdrawer_119,hanger_111]=True
    close[closetdrawer_119,hanger_112]=True
    close[closetdrawer_119,hanger_113]=True
    close[closetdrawer_119,hanger_114]=True
    close[closetdrawer_119,hanger_115]=True
    close[closetdrawer_119,closetdrawer_116]=True
    close[closetdrawer_119,closetdrawer_117]=True
    close[closetdrawer_119,closetdrawer_118]=True
    close[closetdrawer_119,closetdrawer_120]=True
    close[closetdrawer_119,closetdrawer_121]=True
    close[closetdrawer_119,closetdrawer_122]=True
    close[closetdrawer_119,dresser_123]=True
    close[closetdrawer_119,hanger_126]=True
    close[closetdrawer_119,hanger_130]=True
    close[closetdrawer_119,hanger_132]=True
    close[closetdrawer_119,hanger_134]=True
    close[closetdrawer_119,hanger_136]=True
    close[closetdrawer_119,closetdrawer_143]=True
    close[closetdrawer_119,closetdrawer_150]=True
    close[closetdrawer_119,closetdrawer_154]=True
    close[closetdrawer_119,closetdrawer_160]=True
    close[closetdrawer_120,floor_68]=True
    close[closetdrawer_120,floor_69]=True
    close[closetdrawer_120,floor_74]=True
    close[closetdrawer_120,wall_78]=True
    close[closetdrawer_120,wall_81]=True
    close[closetdrawer_120,dresser_108]=True
    close[closetdrawer_120,hanger_109]=True
    close[closetdrawer_120,hanger_110]=True
    close[closetdrawer_120,hanger_111]=True
    close[closetdrawer_120,hanger_112]=True
    close[closetdrawer_120,hanger_113]=True
    close[closetdrawer_120,hanger_114]=True
    close[closetdrawer_120,hanger_115]=True
    close[closetdrawer_120,closetdrawer_116]=True
    close[closetdrawer_120,closetdrawer_117]=True
    close[closetdrawer_120,closetdrawer_118]=True
    close[closetdrawer_120,closetdrawer_119]=True
    close[closetdrawer_120,closetdrawer_121]=True
    close[closetdrawer_120,closetdrawer_122]=True
    close[closetdrawer_120,dresser_123]=True
    close[closetdrawer_120,hanger_132]=True
    close[closetdrawer_120,closetdrawer_143]=True
    close[closetdrawer_120,closetdrawer_150]=True
    close[closetdrawer_120,closetdrawer_154]=True
    close[closetdrawer_120,closetdrawer_160]=True
    close[closetdrawer_121,floor_68]=True
    close[closetdrawer_121,floor_69]=True
    close[closetdrawer_121,floor_74]=True
    close[closetdrawer_121,wall_78]=True
    close[closetdrawer_121,wall_81]=True
    close[closetdrawer_121,dresser_108]=True
    close[closetdrawer_121,closetdrawer_116]=True
    close[closetdrawer_121,closetdrawer_117]=True
    close[closetdrawer_121,closetdrawer_118]=True
    close[closetdrawer_121,closetdrawer_119]=True
    close[closetdrawer_121,closetdrawer_120]=True
    close[closetdrawer_121,closetdrawer_122]=True
    close[closetdrawer_121,dresser_123]=True
    close[closetdrawer_121,closetdrawer_143]=True
    close[closetdrawer_121,closetdrawer_146]=True
    close[closetdrawer_121,closetdrawer_148]=True
    close[closetdrawer_121,closetdrawer_150]=True
    close[closetdrawer_121,closetdrawer_154]=True
    close[closetdrawer_121,closetdrawer_158]=True
    close[closetdrawer_121,closetdrawer_160]=True
    close[closetdrawer_121,mat_173]=True
    close[closetdrawer_122,floor_68]=True
    close[closetdrawer_122,floor_69]=True
    close[closetdrawer_122,floor_74]=True
    close[closetdrawer_122,wall_78]=True
    close[closetdrawer_122,wall_81]=True
    close[closetdrawer_122,dresser_108]=True
    close[closetdrawer_122,closetdrawer_116]=True
    close[closetdrawer_122,closetdrawer_117]=True
    close[closetdrawer_122,closetdrawer_118]=True
    close[closetdrawer_122,closetdrawer_119]=True
    close[closetdrawer_122,closetdrawer_120]=True
    close[closetdrawer_122,closetdrawer_121]=True
    close[closetdrawer_122,dresser_123]=True
    close[closetdrawer_122,closetdrawer_143]=True
    close[closetdrawer_122,closetdrawer_150]=True
    close[closetdrawer_122,closetdrawer_154]=True
    close[closetdrawer_122,closetdrawer_160]=True
    close[closetdrawer_122,mat_173]=True
    close[dresser_123,floor_68]=True
    close[dresser_123,floor_69]=True
    close[dresser_123,wall_81]=True
    close[dresser_123,ceiling_87]=True
    close[dresser_123,dresser_108]=True
    close[dresser_123,hanger_109]=True
    close[dresser_123,hanger_110]=True
    close[dresser_123,hanger_111]=True
    close[dresser_123,hanger_112]=True
    close[dresser_123,hanger_113]=True
    close[dresser_123,hanger_114]=True
    close[dresser_123,hanger_115]=True
    close[dresser_123,closetdrawer_116]=True
    close[dresser_123,closetdrawer_117]=True
    close[dresser_123,closetdrawer_118]=True
    close[dresser_123,closetdrawer_119]=True
    close[dresser_123,closetdrawer_120]=True
    close[dresser_123,closetdrawer_121]=True
    close[dresser_123,closetdrawer_122]=True
    close[dresser_123,hanger_124]=True
    close[dresser_123,hanger_126]=True
    close[dresser_123,hanger_128]=True
    close[dresser_123,hanger_130]=True
    close[dresser_123,hanger_132]=True
    close[dresser_123,hanger_134]=True
    close[dresser_123,hanger_136]=True
    close[dresser_123,hanger_138]=True
    close[dresser_123,hanger_140]=True
    close[dresser_123,hanger_141]=True
    close[dresser_123,hanger_142]=True
    close[dresser_123,closetdrawer_143]=True
    close[dresser_123,closetdrawer_146]=True
    close[dresser_123,closetdrawer_148]=True
    close[dresser_123,closetdrawer_150]=True
    close[dresser_123,closetdrawer_154]=True
    close[dresser_123,closetdrawer_158]=True
    close[dresser_123,closetdrawer_160]=True
    close[hanger_124,wall_81]=True
    close[hanger_124,ceiling_87]=True
    close[hanger_124,dresser_108]=True
    close[hanger_124,closetdrawer_117]=True
    close[hanger_124,dresser_123]=True
    close[hanger_124,hanger_126]=True
    close[hanger_124,hanger_128]=True
    close[hanger_124,hanger_130]=True
    close[hanger_124,hanger_132]=True
    close[hanger_124,hanger_134]=True
    close[hanger_124,hanger_136]=True
    close[hanger_124,hanger_138]=True
    close[hanger_124,hanger_140]=True
    close[hanger_124,hanger_141]=True
    close[hanger_124,hanger_142]=True
    close[hanger_124,closetdrawer_143]=True
    close[hanger_124,closetdrawer_146]=True
    close[hanger_124,closetdrawer_148]=True
    close[hanger_124,closetdrawer_150]=True
    close[hanger_124,closetdrawer_154]=True
    close[hanger_126,wall_78]=True
    close[hanger_126,wall_81]=True
    close[hanger_126,ceiling_87]=True
    close[hanger_126,ceiling_92]=True
    close[hanger_126,dresser_108]=True
    close[hanger_126,hanger_109]=True
    close[hanger_126,hanger_110]=True
    close[hanger_126,hanger_111]=True
    close[hanger_126,hanger_112]=True
    close[hanger_126,hanger_113]=True
    close[hanger_126,hanger_115]=True
    close[hanger_126,closetdrawer_116]=True
    close[hanger_126,closetdrawer_117]=True
    close[hanger_126,closetdrawer_118]=True
    close[hanger_126,closetdrawer_119]=True
    close[hanger_126,dresser_123]=True
    close[hanger_126,hanger_124]=True
    close[hanger_126,hanger_128]=True
    close[hanger_126,hanger_130]=True
    close[hanger_126,hanger_132]=True
    close[hanger_126,hanger_134]=True
    close[hanger_126,hanger_136]=True
    close[hanger_126,hanger_138]=True
    close[hanger_126,hanger_140]=True
    close[hanger_126,hanger_141]=True
    close[hanger_126,hanger_142]=True
    close[hanger_126,closetdrawer_143]=True
    close[hanger_126,closetdrawer_146]=True
    close[hanger_126,closetdrawer_150]=True
    close[hanger_126,closetdrawer_154]=True
    close[hanger_128,wall_81]=True
    close[hanger_128,ceiling_87]=True
    close[hanger_128,dresser_108]=True
    close[hanger_128,hanger_109]=True
    close[hanger_128,hanger_110]=True
    close[hanger_128,closetdrawer_117]=True
    close[hanger_128,dresser_123]=True
    close[hanger_128,hanger_124]=True
    close[hanger_128,hanger_126]=True
    close[hanger_128,hanger_130]=True
    close[hanger_128,hanger_132]=True
    close[hanger_128,hanger_134]=True
    close[hanger_128,hanger_136]=True
    close[hanger_128,hanger_138]=True
    close[hanger_128,hanger_140]=True
    close[hanger_128,hanger_141]=True
    close[hanger_128,hanger_142]=True
    close[hanger_128,closetdrawer_143]=True
    close[hanger_128,closetdrawer_146]=True
    close[hanger_128,closetdrawer_148]=True
    close[hanger_128,closetdrawer_150]=True
    close[hanger_128,closetdrawer_154]=True
    close[hanger_130,wall_78]=True
    close[hanger_130,wall_81]=True
    close[hanger_130,ceiling_87]=True
    close[hanger_130,ceiling_92]=True
    close[hanger_130,dresser_108]=True
    close[hanger_130,hanger_109]=True
    close[hanger_130,hanger_110]=True
    close[hanger_130,hanger_111]=True
    close[hanger_130,hanger_112]=True
    close[hanger_130,hanger_113]=True
    close[hanger_130,closetdrawer_116]=True
    close[hanger_130,closetdrawer_117]=True
    close[hanger_130,closetdrawer_118]=True
    close[hanger_130,closetdrawer_119]=True
    close[hanger_130,dresser_123]=True
    close[hanger_130,hanger_124]=True
    close[hanger_130,hanger_126]=True
    close[hanger_130,hanger_128]=True
    close[hanger_130,hanger_132]=True
    close[hanger_130,hanger_134]=True
    close[hanger_130,hanger_136]=True
    close[hanger_130,hanger_138]=True
    close[hanger_130,hanger_140]=True
    close[hanger_130,hanger_141]=True
    close[hanger_130,hanger_142]=True
    close[hanger_130,closetdrawer_143]=True
    close[hanger_130,closetdrawer_146]=True
    close[hanger_130,closetdrawer_148]=True
    close[hanger_130,closetdrawer_150]=True
    close[hanger_130,closetdrawer_154]=True
    close[hanger_132,wall_78]=True
    close[hanger_132,wall_81]=True
    close[hanger_132,ceiling_87]=True
    close[hanger_132,ceiling_92]=True
    close[hanger_132,dresser_108]=True
    close[hanger_132,hanger_109]=True
    close[hanger_132,hanger_110]=True
    close[hanger_132,hanger_111]=True
    close[hanger_132,hanger_112]=True
    close[hanger_132,hanger_113]=True
    close[hanger_132,hanger_114]=True
    close[hanger_132,hanger_115]=True
    close[hanger_132,closetdrawer_116]=True
    close[hanger_132,closetdrawer_117]=True
    close[hanger_132,closetdrawer_118]=True
    close[hanger_132,closetdrawer_119]=True
    close[hanger_132,closetdrawer_120]=True
    close[hanger_132,dresser_123]=True
    close[hanger_132,hanger_124]=True
    close[hanger_132,hanger_126]=True
    close[hanger_132,hanger_128]=True
    close[hanger_132,hanger_130]=True
    close[hanger_132,hanger_134]=True
    close[hanger_132,hanger_136]=True
    close[hanger_132,hanger_138]=True
    close[hanger_132,hanger_140]=True
    close[hanger_132,hanger_141]=True
    close[hanger_132,hanger_142]=True
    close[hanger_132,closetdrawer_143]=True
    close[hanger_132,closetdrawer_146]=True
    close[hanger_132,closetdrawer_150]=True
    close[hanger_132,closetdrawer_154]=True
    close[hanger_134,wall_78]=True
    close[hanger_134,wall_81]=True
    close[hanger_134,ceiling_87]=True
    close[hanger_134,ceiling_92]=True
    close[hanger_134,dresser_108]=True
    close[hanger_134,hanger_109]=True
    close[hanger_134,hanger_110]=True
    close[hanger_134,hanger_111]=True
    close[hanger_134,hanger_112]=True
    close[hanger_134,hanger_113]=True
    close[hanger_134,hanger_115]=True
    close[hanger_134,closetdrawer_116]=True
    close[hanger_134,closetdrawer_117]=True
    close[hanger_134,closetdrawer_118]=True
    close[hanger_134,closetdrawer_119]=True
    close[hanger_134,dresser_123]=True
    close[hanger_134,hanger_124]=True
    close[hanger_134,hanger_126]=True
    close[hanger_134,hanger_128]=True
    close[hanger_134,hanger_130]=True
    close[hanger_134,hanger_132]=True
    close[hanger_134,hanger_136]=True
    close[hanger_134,hanger_138]=True
    close[hanger_134,hanger_140]=True
    close[hanger_134,hanger_141]=True
    close[hanger_134,hanger_142]=True
    close[hanger_134,closetdrawer_143]=True
    close[hanger_134,closetdrawer_146]=True
    close[hanger_134,closetdrawer_150]=True
    close[hanger_134,closetdrawer_154]=True
    close[hanger_136,wall_78]=True
    close[hanger_136,wall_81]=True
    close[hanger_136,ceiling_87]=True
    close[hanger_136,dresser_108]=True
    close[hanger_136,hanger_109]=True
    close[hanger_136,hanger_110]=True
    close[hanger_136,hanger_111]=True
    close[hanger_136,hanger_112]=True
    close[hanger_136,closetdrawer_116]=True
    close[hanger_136,closetdrawer_117]=True
    close[hanger_136,closetdrawer_118]=True
    close[hanger_136,closetdrawer_119]=True
    close[hanger_136,dresser_123]=True
    close[hanger_136,hanger_124]=True
    close[hanger_136,hanger_126]=True
    close[hanger_136,hanger_128]=True
    close[hanger_136,hanger_130]=True
    close[hanger_136,hanger_132]=True
    close[hanger_136,hanger_134]=True
    close[hanger_136,hanger_138]=True
    close[hanger_136,hanger_140]=True
    close[hanger_136,hanger_141]=True
    close[hanger_136,hanger_142]=True
    close[hanger_136,closetdrawer_143]=True
    close[hanger_136,closetdrawer_146]=True
    close[hanger_136,closetdrawer_148]=True
    close[hanger_136,closetdrawer_150]=True
    close[hanger_136,closetdrawer_154]=True
    close[hanger_138,wall_81]=True
    close[hanger_138,ceiling_87]=True
    close[hanger_138,dresser_108]=True
    close[hanger_138,hanger_109]=True
    close[hanger_138,hanger_110]=True
    close[hanger_138,hanger_111]=True
    close[hanger_138,closetdrawer_116]=True
    close[hanger_138,closetdrawer_117]=True
    close[hanger_138,closetdrawer_118]=True
    close[hanger_138,dresser_123]=True
    close[hanger_138,hanger_124]=True
    close[hanger_138,hanger_126]=True
    close[hanger_138,hanger_128]=True
    close[hanger_138,hanger_130]=True
    close[hanger_138,hanger_132]=True
    close[hanger_138,hanger_134]=True
    close[hanger_138,hanger_136]=True
    close[hanger_138,hanger_140]=True
    close[hanger_138,hanger_141]=True
    close[hanger_138,hanger_142]=True
    close[hanger_138,closetdrawer_143]=True
    close[hanger_138,closetdrawer_146]=True
    close[hanger_138,closetdrawer_148]=True
    close[hanger_138,closetdrawer_150]=True
    close[hanger_138,closetdrawer_154]=True
    close[hanger_140,wall_81]=True
    close[hanger_140,ceiling_87]=True
    close[hanger_140,dresser_108]=True
    close[hanger_140,dresser_123]=True
    close[hanger_140,hanger_124]=True
    close[hanger_140,hanger_126]=True
    close[hanger_140,hanger_128]=True
    close[hanger_140,hanger_130]=True
    close[hanger_140,hanger_132]=True
    close[hanger_140,hanger_134]=True
    close[hanger_140,hanger_136]=True
    close[hanger_140,hanger_138]=True
    close[hanger_140,hanger_141]=True
    close[hanger_140,hanger_142]=True
    close[hanger_140,closetdrawer_143]=True
    close[hanger_140,closetdrawer_146]=True
    close[hanger_140,closetdrawer_148]=True
    close[hanger_140,closetdrawer_150]=True
    close[hanger_140,closetdrawer_154]=True
    close[hanger_141,wall_81]=True
    close[hanger_141,ceiling_87]=True
    close[hanger_141,dresser_108]=True
    close[hanger_141,dresser_123]=True
    close[hanger_141,hanger_124]=True
    close[hanger_141,hanger_126]=True
    close[hanger_141,hanger_128]=True
    close[hanger_141,hanger_130]=True
    close[hanger_141,hanger_132]=True
    close[hanger_141,hanger_134]=True
    close[hanger_141,hanger_136]=True
    close[hanger_141,hanger_138]=True
    close[hanger_141,hanger_140]=True
    close[hanger_141,hanger_142]=True
    close[hanger_141,closetdrawer_143]=True
    close[hanger_141,closetdrawer_146]=True
    close[hanger_141,closetdrawer_148]=True
    close[hanger_141,closetdrawer_150]=True
    close[hanger_141,closetdrawer_154]=True
    close[hanger_142,wall_81]=True
    close[hanger_142,ceiling_87]=True
    close[hanger_142,dresser_108]=True
    close[hanger_142,dresser_123]=True
    close[hanger_142,hanger_124]=True
    close[hanger_142,hanger_126]=True
    close[hanger_142,hanger_128]=True
    close[hanger_142,hanger_130]=True
    close[hanger_142,hanger_132]=True
    close[hanger_142,hanger_134]=True
    close[hanger_142,hanger_136]=True
    close[hanger_142,hanger_138]=True
    close[hanger_142,hanger_140]=True
    close[hanger_142,hanger_141]=True
    close[hanger_142,closetdrawer_143]=True
    close[hanger_142,closetdrawer_146]=True
    close[hanger_142,closetdrawer_148]=True
    close[hanger_142,closetdrawer_150]=True
    close[hanger_142,closetdrawer_154]=True
    close[closetdrawer_143,floor_68]=True
    close[closetdrawer_143,floor_69]=True
    close[closetdrawer_143,wall_78]=True
    close[closetdrawer_143,wall_81]=True
    close[closetdrawer_143,dresser_108]=True
    close[closetdrawer_143,hanger_109]=True
    close[closetdrawer_143,hanger_110]=True
    close[closetdrawer_143,hanger_111]=True
    close[closetdrawer_143,hanger_112]=True
    close[closetdrawer_143,hanger_113]=True
    close[closetdrawer_143,closetdrawer_116]=True
    close[closetdrawer_143,closetdrawer_117]=True
    close[closetdrawer_143,closetdrawer_118]=True
    close[closetdrawer_143,closetdrawer_119]=True
    close[closetdrawer_143,closetdrawer_120]=True
    close[closetdrawer_143,closetdrawer_121]=True
    close[closetdrawer_143,closetdrawer_122]=True
    close[closetdrawer_143,dresser_123]=True
    close[closetdrawer_143,hanger_124]=True
    close[closetdrawer_143,hanger_126]=True
    close[closetdrawer_143,hanger_128]=True
    close[closetdrawer_143,hanger_130]=True
    close[closetdrawer_143,hanger_132]=True
    close[closetdrawer_143,hanger_134]=True
    close[closetdrawer_143,hanger_136]=True
    close[closetdrawer_143,hanger_138]=True
    close[closetdrawer_143,hanger_140]=True
    close[closetdrawer_143,hanger_141]=True
    close[closetdrawer_143,hanger_142]=True
    close[closetdrawer_143,closetdrawer_146]=True
    close[closetdrawer_143,closetdrawer_148]=True
    close[closetdrawer_143,closetdrawer_150]=True
    close[closetdrawer_143,closetdrawer_154]=True
    close[closetdrawer_143,closetdrawer_158]=True
    close[closetdrawer_143,closetdrawer_160]=True
    close[closetdrawer_146,floor_68]=True
    close[closetdrawer_146,floor_69]=True
    close[closetdrawer_146,wall_81]=True
    close[closetdrawer_146,dresser_108]=True
    close[closetdrawer_146,closetdrawer_117]=True
    close[closetdrawer_146,closetdrawer_118]=True
    close[closetdrawer_146,closetdrawer_121]=True
    close[closetdrawer_146,dresser_123]=True
    close[closetdrawer_146,hanger_124]=True
    close[closetdrawer_146,hanger_126]=True
    close[closetdrawer_146,hanger_128]=True
    close[closetdrawer_146,hanger_130]=True
    close[closetdrawer_146,hanger_132]=True
    close[closetdrawer_146,hanger_134]=True
    close[closetdrawer_146,hanger_136]=True
    close[closetdrawer_146,hanger_138]=True
    close[closetdrawer_146,hanger_140]=True
    close[closetdrawer_146,hanger_141]=True
    close[closetdrawer_146,hanger_142]=True
    close[closetdrawer_146,closetdrawer_143]=True
    close[closetdrawer_146,closetdrawer_148]=True
    close[closetdrawer_146,closetdrawer_150]=True
    close[closetdrawer_146,closetdrawer_154]=True
    close[closetdrawer_146,closetdrawer_158]=True
    close[closetdrawer_146,closetdrawer_160]=True
    close[closetdrawer_148,floor_68]=True
    close[closetdrawer_148,floor_69]=True
    close[closetdrawer_148,wall_81]=True
    close[closetdrawer_148,dresser_108]=True
    close[closetdrawer_148,closetdrawer_117]=True
    close[closetdrawer_148,closetdrawer_118]=True
    close[closetdrawer_148,closetdrawer_121]=True
    close[closetdrawer_148,dresser_123]=True
    close[closetdrawer_148,hanger_124]=True
    close[closetdrawer_148,hanger_128]=True
    close[closetdrawer_148,hanger_130]=True
    close[closetdrawer_148,hanger_136]=True
    close[closetdrawer_148,hanger_138]=True
    close[closetdrawer_148,hanger_140]=True
    close[closetdrawer_148,hanger_141]=True
    close[closetdrawer_148,hanger_142]=True
    close[closetdrawer_148,closetdrawer_143]=True
    close[closetdrawer_148,closetdrawer_146]=True
    close[closetdrawer_148,closetdrawer_150]=True
    close[closetdrawer_148,closetdrawer_154]=True
    close[closetdrawer_148,closetdrawer_158]=True
    close[closetdrawer_148,closetdrawer_160]=True
    close[closetdrawer_150,floor_68]=True
    close[closetdrawer_150,floor_69]=True
    close[closetdrawer_150,wall_78]=True
    close[closetdrawer_150,wall_81]=True
    close[closetdrawer_150,dresser_108]=True
    close[closetdrawer_150,hanger_109]=True
    close[closetdrawer_150,hanger_110]=True
    close[closetdrawer_150,hanger_111]=True
    close[closetdrawer_150,hanger_112]=True
    close[closetdrawer_150,closetdrawer_116]=True
    close[closetdrawer_150,closetdrawer_117]=True
    close[closetdrawer_150,closetdrawer_118]=True
    close[closetdrawer_150,closetdrawer_119]=True
    close[closetdrawer_150,closetdrawer_120]=True
    close[closetdrawer_150,closetdrawer_121]=True
    close[closetdrawer_150,closetdrawer_122]=True
    close[closetdrawer_150,dresser_123]=True
    close[closetdrawer_150,hanger_124]=True
    close[closetdrawer_150,hanger_126]=True
    close[closetdrawer_150,hanger_128]=True
    close[closetdrawer_150,hanger_130]=True
    close[closetdrawer_150,hanger_132]=True
    close[closetdrawer_150,hanger_134]=True
    close[closetdrawer_150,hanger_136]=True
    close[closetdrawer_150,hanger_138]=True
    close[closetdrawer_150,hanger_140]=True
    close[closetdrawer_150,hanger_141]=True
    close[closetdrawer_150,hanger_142]=True
    close[closetdrawer_150,closetdrawer_143]=True
    close[closetdrawer_150,closetdrawer_146]=True
    close[closetdrawer_150,closetdrawer_148]=True
    close[closetdrawer_150,closetdrawer_154]=True
    close[closetdrawer_150,closetdrawer_158]=True
    close[closetdrawer_150,closetdrawer_160]=True
    close[closetdrawer_154,floor_68]=True
    close[closetdrawer_154,floor_69]=True
    close[closetdrawer_154,floor_74]=True
    close[closetdrawer_154,wall_78]=True
    close[closetdrawer_154,wall_81]=True
    close[closetdrawer_154,dresser_108]=True
    close[closetdrawer_154,hanger_109]=True
    close[closetdrawer_154,closetdrawer_116]=True
    close[closetdrawer_154,closetdrawer_117]=True
    close[closetdrawer_154,closetdrawer_118]=True
    close[closetdrawer_154,closetdrawer_119]=True
    close[closetdrawer_154,closetdrawer_120]=True
    close[closetdrawer_154,closetdrawer_121]=True
    close[closetdrawer_154,closetdrawer_122]=True
    close[closetdrawer_154,dresser_123]=True
    close[closetdrawer_154,hanger_124]=True
    close[closetdrawer_154,hanger_126]=True
    close[closetdrawer_154,hanger_128]=True
    close[closetdrawer_154,hanger_130]=True
    close[closetdrawer_154,hanger_132]=True
    close[closetdrawer_154,hanger_134]=True
    close[closetdrawer_154,hanger_136]=True
    close[closetdrawer_154,hanger_138]=True
    close[closetdrawer_154,hanger_140]=True
    close[closetdrawer_154,hanger_141]=True
    close[closetdrawer_154,hanger_142]=True
    close[closetdrawer_154,closetdrawer_143]=True
    close[closetdrawer_154,closetdrawer_146]=True
    close[closetdrawer_154,closetdrawer_148]=True
    close[closetdrawer_154,closetdrawer_150]=True
    close[closetdrawer_154,closetdrawer_158]=True
    close[closetdrawer_154,closetdrawer_160]=True
    close[closetdrawer_158,floor_68]=True
    close[closetdrawer_158,floor_69]=True
    close[closetdrawer_158,wall_81]=True
    close[closetdrawer_158,dresser_108]=True
    close[closetdrawer_158,closetdrawer_117]=True
    close[closetdrawer_158,closetdrawer_118]=True
    close[closetdrawer_158,closetdrawer_121]=True
    close[closetdrawer_158,dresser_123]=True
    close[closetdrawer_158,closetdrawer_143]=True
    close[closetdrawer_158,closetdrawer_146]=True
    close[closetdrawer_158,closetdrawer_148]=True
    close[closetdrawer_158,closetdrawer_150]=True
    close[closetdrawer_158,closetdrawer_154]=True
    close[closetdrawer_158,closetdrawer_160]=True
    close[closetdrawer_158,mat_173]=True
    close[closetdrawer_160,floor_68]=True
    close[closetdrawer_160,floor_69]=True
    close[closetdrawer_160,floor_74]=True
    close[closetdrawer_160,wall_78]=True
    close[closetdrawer_160,wall_81]=True
    close[closetdrawer_160,dresser_108]=True
    close[closetdrawer_160,closetdrawer_116]=True
    close[closetdrawer_160,closetdrawer_117]=True
    close[closetdrawer_160,closetdrawer_118]=True
    close[closetdrawer_160,closetdrawer_119]=True
    close[closetdrawer_160,closetdrawer_120]=True
    close[closetdrawer_160,closetdrawer_121]=True
    close[closetdrawer_160,closetdrawer_122]=True
    close[closetdrawer_160,dresser_123]=True
    close[closetdrawer_160,closetdrawer_143]=True
    close[closetdrawer_160,closetdrawer_146]=True
    close[closetdrawer_160,closetdrawer_148]=True
    close[closetdrawer_160,closetdrawer_150]=True
    close[closetdrawer_160,closetdrawer_154]=True
    close[closetdrawer_160,closetdrawer_158]=True
    close[closetdrawer_160,mat_173]=True
    close[doorjamb_165,floor_76]=True
    close[doorjamb_165,wall_83]=True
    close[doorjamb_165,wall_84]=True
    close[doorjamb_165,wall_85]=True
    close[doorjamb_165,ceiling_94]=True
    close[doorjamb_165,trashcan_99]=True
    close[doorjamb_165,desk_104]=True
    close[doorjamb_165,light_169]=True
    close[doorjamb_165,computer_170]=True
    close[doorjamb_165,drawing_174]=True
    close[doorjamb_165,floor_206]=True
    close[doorjamb_165,wall_209]=True
    close[doorjamb_165,wall_210]=True
    close[doorjamb_165,wall_211]=True
    close[doorjamb_165,ceiling_217]=True
    close[doorjamb_165,door_222]=True
    close[doorjamb_165,bookshelf_233]=True
    close[doorjamb_165,drawing_238]=True
    close[doorjamb_165,drawing_240]=True
    close[doorjamb_165,light_245]=True
    close[doorjamb_165,powersocket_246]=True
    close[doorjamb_165,phone_247]=True
    close[doorjamb_165,wall_clock_249]=True
    close[mouse_166,floor_75]=True
    close[mouse_166,wall_83]=True
    close[mouse_166,chair_103]=True
    close[mouse_166,desk_104]=True
    close[mouse_166,mousepad_167]=True
    close[mouse_166,keyboard_168]=True
    close[mouse_166,computer_170]=True
    close[mouse_166,cpuscreen_171]=True
    close[mouse_166,drawing_175]=True
    close[mouse_166,floor_207]=True
    close[mouse_166,wall_210]=True
    close[mouse_166,bookshelf_233]=True
    close[mousepad_167,floor_75]=True
    close[mousepad_167,wall_83]=True
    close[mousepad_167,chair_103]=True
    close[mousepad_167,desk_104]=True
    close[mousepad_167,mouse_166]=True
    close[mousepad_167,keyboard_168]=True
    close[mousepad_167,computer_170]=True
    close[mousepad_167,cpuscreen_171]=True
    close[mousepad_167,drawing_175]=True
    close[mousepad_167,floor_207]=True
    close[mousepad_167,wall_210]=True
    close[mousepad_167,bookshelf_233]=True
    close[keyboard_168,floor_75]=True
    close[keyboard_168,floor_76]=True
    close[keyboard_168,wall_83]=True
    close[keyboard_168,wall_84]=True
    close[keyboard_168,chair_103]=True
    close[keyboard_168,desk_104]=True
    close[keyboard_168,mouse_166]=True
    close[keyboard_168,mousepad_167]=True
    close[keyboard_168,light_169]=True
    close[keyboard_168,computer_170]=True
    close[keyboard_168,cpuscreen_171]=True
    close[keyboard_168,floor_207]=True
    close[keyboard_168,wall_209]=True
    close[keyboard_168,wall_210]=True
    close[keyboard_168,bookshelf_233]=True
    close[light_169,floor_75]=True
    close[light_169,floor_76]=True
    close[light_169,wall_83]=True
    close[light_169,wall_84]=True
    close[light_169,ceiling_93]=True
    close[light_169,ceiling_94]=True
    close[light_169,chair_103]=True
    close[light_169,desk_104]=True
    close[light_169,doorjamb_165]=True
    close[light_169,keyboard_168]=True
    close[light_169,computer_170]=True
    close[light_169,cpuscreen_171]=True
    close[light_169,drawing_174]=True
    close[light_169,floor_206]=True
    close[light_169,floor_207]=True
    close[light_169,wall_209]=True
    close[light_169,wall_210]=True
    close[light_169,ceiling_217]=True
    close[light_169,ceiling_218]=True
    close[light_169,door_222]=True
    close[light_169,bookshelf_233]=True
    close[light_169,light_245]=True
    close[light_169,powersocket_246]=True
    close[light_169,phone_247]=True
    close[computer_170,floor_75]=True
    close[computer_170,floor_76]=True
    close[computer_170,wall_83]=True
    close[computer_170,wall_84]=True
    close[computer_170,chair_103]=True
    close[computer_170,desk_104]=True
    close[computer_170,doorjamb_165]=True
    close[computer_170,mouse_166]=True
    close[computer_170,mousepad_167]=True
    close[computer_170,keyboard_168]=True
    close[computer_170,light_169]=True
    close[computer_170,cpuscreen_171]=True
    close[computer_170,floor_206]=True
    close[computer_170,floor_207]=True
    close[computer_170,wall_209]=True
    close[computer_170,wall_210]=True
    close[computer_170,door_222]=True
    close[computer_170,bookshelf_233]=True
    close[cpuscreen_171,floor_75]=True
    close[cpuscreen_171,floor_76]=True
    close[cpuscreen_171,wall_83]=True
    close[cpuscreen_171,wall_84]=True
    close[cpuscreen_171,ceiling_93]=True
    close[cpuscreen_171,chair_103]=True
    close[cpuscreen_171,desk_104]=True
    close[cpuscreen_171,mouse_166]=True
    close[cpuscreen_171,mousepad_167]=True
    close[cpuscreen_171,keyboard_168]=True
    close[cpuscreen_171,light_169]=True
    close[cpuscreen_171,computer_170]=True
    close[cpuscreen_171,floor_207]=True
    close[cpuscreen_171,wall_209]=True
    close[cpuscreen_171,wall_210]=True
    close[cpuscreen_171,ceiling_218]=True
    close[cpuscreen_171,bookshelf_233]=True
    close[mat_173,floor_68]=True
    close[mat_173,floor_69]=True
    close[mat_173,floor_70]=True
    close[mat_173,floor_71]=True
    close[mat_173,floor_72]=True
    close[mat_173,floor_73]=True
    close[mat_173,floor_74]=True
    close[mat_173,wall_80]=True
    close[mat_173,wall_81]=True
    close[mat_173,wall_82]=True
    close[mat_173,window_86]=True
    close[mat_173,tablelamp_97]=True
    close[mat_173,tablelamp_98]=True
    close[mat_173,nightstand_100]=True
    close[mat_173,nightstand_102]=True
    close[mat_173,bed_105]=True
    close[mat_173,chair_106]=True
    close[mat_173,table_107]=True
    close[mat_173,closetdrawer_121]=True
    close[mat_173,closetdrawer_122]=True
    close[mat_173,closetdrawer_158]=True
    close[mat_173,closetdrawer_160]=True
    close[mat_173,orchid_178]=True
    close[mat_173,curtain_179]=True
    close[mat_173,curtain_180]=True
    close[mat_173,curtain_181]=True
    close[mat_173,pillow_182]=True
    close[mat_173,pillow_183]=True
    close[drawing_174,wall_14]=True
    close[drawing_174,door_44]=True
    close[drawing_174,doorjamb_45]=True
    close[drawing_174,floor_76]=True
    close[drawing_174,floor_77]=True
    close[drawing_174,wall_84]=True
    close[drawing_174,wall_85]=True
    close[drawing_174,ceiling_94]=True
    close[drawing_174,ceiling_95]=True
    close[drawing_174,trashcan_99]=True
    close[drawing_174,doorjamb_165]=True
    close[drawing_174,light_169]=True
    close[drawing_174,floor_202]=True
    close[drawing_174,floor_203]=True
    close[drawing_174,floor_206]=True
    close[drawing_174,wall_209]=True
    close[drawing_174,wall_211]=True
    close[drawing_174,ceiling_216]=True
    close[drawing_174,ceiling_217]=True
    close[drawing_174,door_222]=True
    close[drawing_174,kitchen_counter_230]=True
    close[drawing_174,drawing_238]=True
    close[drawing_174,drawing_239]=True
    close[drawing_174,drawing_240]=True
    close[drawing_174,light_245]=True
    close[drawing_174,powersocket_246]=True
    close[drawing_174,phone_247]=True
    close[drawing_174,wall_clock_249]=True
    close[drawing_174,fridge_289]=True
    close[drawing_174,microwave_297]=True
    close[drawing_175,floor_74]=True
    close[drawing_175,floor_75]=True
    close[drawing_175,wall_78]=True
    close[drawing_175,wall_83]=True
    close[drawing_175,ceiling_92]=True
    close[drawing_175,ceiling_93]=True
    close[drawing_175,desk_104]=True
    close[drawing_175,mouse_166]=True
    close[drawing_175,mousepad_167]=True
    close[drawing_176,floor_2]=True
    close[drawing_176,floor_3]=True
    close[drawing_176,wall_12]=True
    close[drawing_176,ceiling_16]=True
    close[drawing_176,walllamp_28]=True
    close[drawing_176,towel_rack_31]=True
    close[drawing_176,bathroom_cabinet_40]=True
    close[drawing_176,bathroom_counter_41]=True
    close[drawing_176,floor_71]=True
    close[drawing_176,wall_79]=True
    close[drawing_176,wall_82]=True
    close[drawing_176,ceiling_89]=True
    close[drawing_176,bookshelf_101]=True
    close[drawing_176,chair_106]=True
    close[drawing_176,photoframe_185]=True
    close[orchid_178,floor_72]=True
    close[orchid_178,floor_73]=True
    close[orchid_178,floor_74]=True
    close[orchid_178,floor_76]=True
    close[orchid_178,table_107]=True
    close[orchid_178,mat_173]=True
    close[curtain_179,floor_70]=True
    close[curtain_179,wall_80]=True
    close[curtain_179,wall_81]=True
    close[curtain_179,window_86]=True
    close[curtain_179,ceiling_87]=True
    close[curtain_179,ceiling_88]=True
    close[curtain_179,tablelamp_97]=True
    close[curtain_179,nightstand_100]=True
    close[curtain_179,bed_105]=True
    close[curtain_179,mat_173]=True
    close[curtain_179,curtain_180]=True
    close[curtain_179,curtain_181]=True
    close[curtain_179,pillow_182]=True
    close[curtain_179,pillow_183]=True
    close[curtain_180,floor_70]=True
    close[curtain_180,wall_80]=True
    close[curtain_180,wall_81]=True
    close[curtain_180,window_86]=True
    close[curtain_180,ceiling_87]=True
    close[curtain_180,ceiling_88]=True
    close[curtain_180,tablelamp_97]=True
    close[curtain_180,nightstand_100]=True
    close[curtain_180,bed_105]=True
    close[curtain_180,mat_173]=True
    close[curtain_180,curtain_179]=True
    close[curtain_180,curtain_181]=True
    close[curtain_180,pillow_182]=True
    close[curtain_180,pillow_183]=True
    close[curtain_181,floor_70]=True
    close[curtain_181,wall_80]=True
    close[curtain_181,wall_82]=True
    close[curtain_181,window_86]=True
    close[curtain_181,ceiling_88]=True
    close[curtain_181,ceiling_89]=True
    close[curtain_181,tablelamp_98]=True
    close[curtain_181,nightstand_102]=True
    close[curtain_181,bed_105]=True
    close[curtain_181,mat_173]=True
    close[curtain_181,curtain_179]=True
    close[curtain_181,curtain_180]=True
    close[curtain_181,pillow_182]=True
    close[curtain_181,pillow_183]=True
    close[pillow_182,floor_70]=True
    close[pillow_182,floor_71]=True
    close[pillow_182,wall_80]=True
    close[pillow_182,wall_82]=True
    close[pillow_182,window_86]=True
    close[pillow_182,tablelamp_97]=True
    close[pillow_182,tablelamp_98]=True
    close[pillow_182,nightstand_100]=True
    close[pillow_182,nightstand_102]=True
    close[pillow_182,bed_105]=True
    close[pillow_182,mat_173]=True
    close[pillow_182,curtain_179]=True
    close[pillow_182,curtain_180]=True
    close[pillow_182,curtain_181]=True
    close[pillow_182,pillow_183]=True
    close[pillow_183,floor_68]=True
    close[pillow_183,floor_69]=True
    close[pillow_183,floor_70]=True
    close[pillow_183,wall_80]=True
    close[pillow_183,wall_81]=True
    close[pillow_183,window_86]=True
    close[pillow_183,tablelamp_97]=True
    close[pillow_183,tablelamp_98]=True
    close[pillow_183,nightstand_100]=True
    close[pillow_183,nightstand_102]=True
    close[pillow_183,bed_105]=True
    close[pillow_183,mat_173]=True
    close[pillow_183,curtain_179]=True
    close[pillow_183,curtain_180]=True
    close[pillow_183,curtain_181]=True
    close[pillow_183,pillow_182]=True
    close[photoframe_185,wall_12]=True
    close[photoframe_185,wall_14]=True
    close[photoframe_185,ceiling_16]=True
    close[photoframe_185,walllamp_28]=True
    close[photoframe_185,towel_rack_31]=True
    close[photoframe_185,towel_rack_32]=True
    close[photoframe_185,wall_79]=True
    close[photoframe_185,wall_82]=True
    close[photoframe_185,wall_85]=True
    close[photoframe_185,ceiling_89]=True
    close[photoframe_185,ceiling_90]=True
    close[photoframe_185,bookshelf_101]=True
    close[photoframe_185,drawing_176]=True
    close[floor_202,floor_7]=True
    close[floor_202,wall_11]=True
    close[floor_202,shower_36]=True
    close[floor_202,toilet_37]=True
    close[floor_202,door_44]=True
    close[floor_202,floor_77]=True
    close[floor_202,wall_85]=True
    close[floor_202,trashcan_99]=True
    close[floor_202,drawing_174]=True
    close[floor_202,floor_203]=True
    close[floor_202,floor_204]=True
    close[floor_202,floor_206]=True
    close[floor_202,wall_211]=True
    close[floor_202,wall_212]=True
    close[floor_202,door_222]=True
    close[floor_202,table_226]=True
    close[floor_202,bench_228]=True
    close[floor_202,kitchen_counter_230]=True
    close[floor_202,sink_231]=True
    close[floor_202,faucet_232]=True
    close[floor_202,mat_237]=True
    close[floor_202,drawing_238]=True
    close[floor_202,drawing_239]=True
    close[floor_202,light_245]=True
    close[floor_202,powersocket_246]=True
    close[floor_202,phone_247]=True
    close[floor_202,fridge_289]=True
    close[floor_202,toaster_292]=True
    close[floor_202,microwave_297]=True
    close[floor_203,floor_7]=True
    close[floor_203,wall_11]=True
    close[floor_203,shower_36]=True
    close[floor_203,toilet_37]=True
    close[floor_203,door_44]=True
    close[floor_203,floor_77]=True
    close[floor_203,wall_85]=True
    close[floor_203,trashcan_99]=True
    close[floor_203,drawing_174]=True
    close[floor_203,floor_202]=True
    close[floor_203,floor_204]=True
    close[floor_203,floor_206]=True
    close[floor_203,wall_211]=True
    close[floor_203,wall_212]=True
    close[floor_203,door_222]=True
    close[floor_203,table_226]=True
    close[floor_203,bench_228]=True
    close[floor_203,kitchen_counter_230]=True
    close[floor_203,sink_231]=True
    close[floor_203,faucet_232]=True
    close[floor_203,mat_237]=True
    close[floor_203,drawing_238]=True
    close[floor_203,drawing_239]=True
    close[floor_203,light_245]=True
    close[floor_203,powersocket_246]=True
    close[floor_203,phone_247]=True
    close[floor_203,fridge_289]=True
    close[floor_203,toaster_292]=True
    close[floor_203,microwave_297]=True
    close[floor_204,wall_15]=True
    close[floor_204,toilet_37]=True
    close[floor_204,floor_202]=True
    close[floor_204,floor_203]=True
    close[floor_204,floor_205]=True
    close[floor_204,wall_211]=True
    close[floor_204,wall_212]=True
    close[floor_204,wall_215]=True
    close[floor_204,table_226]=True
    close[floor_204,bench_228]=True
    close[floor_204,kitchen_counter_230]=True
    close[floor_204,sink_231]=True
    close[floor_204,faucet_232]=True
    close[floor_204,mat_237]=True
    close[floor_204,drawing_243]=True
    close[floor_204,coffe_maker_290]=True
    close[floor_204,toaster_292]=True
    close[floor_204,oven_295]=True
    close[floor_204,tray_296]=True
    close[floor_205,floor_204]=True
    close[floor_205,floor_206]=True
    close[floor_205,floor_208]=True
    close[floor_205,wall_212]=True
    close[floor_205,wall_213]=True
    close[floor_205,wall_214]=True
    close[floor_205,table_226]=True
    close[floor_205,bench_227]=True
    close[floor_205,bench_228]=True
    close[floor_205,mat_236]=True
    close[floor_205,mat_237]=True
    close[floor_205,drawing_242]=True
    close[floor_205,drawing_243]=True
    close[floor_205,floor_320]=True
    close[floor_205,wall_332]=True
    close[floor_205,filing_cabinet_399]=True
    close[floor_205,light_411]=True
    close[floor_206,floor_76]=True
    close[floor_206,wall_84]=True
    close[floor_206,trashcan_99]=True
    close[floor_206,desk_104]=True
    close[floor_206,doorjamb_165]=True
    close[floor_206,light_169]=True
    close[floor_206,computer_170]=True
    close[floor_206,drawing_174]=True
    close[floor_206,floor_202]=True
    close[floor_206,floor_203]=True
    close[floor_206,floor_205]=True
    close[floor_206,floor_207]=True
    close[floor_206,wall_209]=True
    close[floor_206,wall_210]=True
    close[floor_206,wall_211]=True
    close[floor_206,door_222]=True
    close[floor_206,table_226]=True
    close[floor_206,bench_227]=True
    close[floor_206,bench_228]=True
    close[floor_206,bookshelf_233]=True
    close[floor_206,mat_236]=True
    close[floor_206,mat_237]=True
    close[floor_206,drawing_238]=True
    close[floor_206,light_245]=True
    close[floor_206,powersocket_246]=True
    close[floor_206,phone_247]=True
    close[floor_207,floor_75]=True
    close[floor_207,wall_83]=True
    close[floor_207,chair_103]=True
    close[floor_207,desk_104]=True
    close[floor_207,mouse_166]=True
    close[floor_207,mousepad_167]=True
    close[floor_207,keyboard_168]=True
    close[floor_207,light_169]=True
    close[floor_207,computer_170]=True
    close[floor_207,cpuscreen_171]=True
    close[floor_207,floor_206]=True
    close[floor_207,floor_208]=True
    close[floor_207,wall_210]=True
    close[floor_207,wall_213]=True
    close[floor_207,door_222]=True
    close[floor_207,tvstand_225]=True
    close[floor_207,table_226]=True
    close[floor_207,bench_227]=True
    close[floor_207,bookshelf_233]=True
    close[floor_207,mat_237]=True
    close[floor_207,orchid_244]=True
    close[floor_207,television_248]=True
    close[floor_207,photoframe_285]=True
    close[floor_208,floor_205]=True
    close[floor_208,floor_207]=True
    close[floor_208,wall_210]=True
    close[floor_208,wall_213]=True
    close[floor_208,tvstand_225]=True
    close[floor_208,table_226]=True
    close[floor_208,bench_227]=True
    close[floor_208,mat_237]=True
    close[floor_208,orchid_244]=True
    close[floor_208,television_248]=True
    close[floor_208,photoframe_285]=True
    close[floor_208,floor_325]=True
    close[floor_208,wall_331]=True
    close[floor_208,doorjamb_346]=True
    close[floor_208,desk_357]=True
    close[floor_208,filing_cabinet_399]=True
    close[floor_208,light_411]=True
    close[floor_208,powersocket_412]=True
    close[floor_208,mouse_413]=True
    close[floor_208,mousepad_414]=True
    close[floor_208,computer_417]=True
    close[wall_209,floor_76]=True
    close[wall_209,wall_83]=True
    close[wall_209,wall_84]=True
    close[wall_209,wall_85]=True
    close[wall_209,ceiling_94]=True
    close[wall_209,trashcan_99]=True
    close[wall_209,chair_103]=True
    close[wall_209,desk_104]=True
    close[wall_209,doorjamb_165]=True
    close[wall_209,keyboard_168]=True
    close[wall_209,light_169]=True
    close[wall_209,computer_170]=True
    close[wall_209,cpuscreen_171]=True
    close[wall_209,drawing_174]=True
    close[wall_209,floor_206]=True
    close[wall_209,wall_210]=True
    close[wall_209,wall_211]=True
    close[wall_209,ceiling_217]=True
    close[wall_209,door_222]=True
    close[wall_209,bookshelf_233]=True
    close[wall_209,drawing_238]=True
    close[wall_209,drawing_239]=True
    close[wall_209,drawing_240]=True
    close[wall_209,light_245]=True
    close[wall_209,powersocket_246]=True
    close[wall_209,phone_247]=True
    close[wall_209,wall_clock_249]=True
    close[wall_210,floor_75]=True
    close[wall_210,wall_83]=True
    close[wall_210,wall_84]=True
    close[wall_210,ceiling_93]=True
    close[wall_210,chair_103]=True
    close[wall_210,desk_104]=True
    close[wall_210,doorjamb_165]=True
    close[wall_210,mouse_166]=True
    close[wall_210,mousepad_167]=True
    close[wall_210,keyboard_168]=True
    close[wall_210,light_169]=True
    close[wall_210,computer_170]=True
    close[wall_210,cpuscreen_171]=True
    close[wall_210,floor_206]=True
    close[wall_210,floor_207]=True
    close[wall_210,floor_208]=True
    close[wall_210,wall_209]=True
    close[wall_210,wall_213]=True
    close[wall_210,ceiling_217]=True
    close[wall_210,ceiling_218]=True
    close[wall_210,ceiling_219]=True
    close[wall_210,door_222]=True
    close[wall_210,ceilinglamp_223]=True
    close[wall_210,tvstand_225]=True
    close[wall_210,table_226]=True
    close[wall_210,bench_227]=True
    close[wall_210,bookshelf_233]=True
    close[wall_210,mat_236]=True
    close[wall_210,mat_237]=True
    close[wall_210,orchid_244]=True
    close[wall_210,television_248]=True
    close[wall_210,photoframe_285]=True
    close[wall_211,floor_7]=True
    close[wall_211,wall_11]=True
    close[wall_211,wall_14]=True
    close[wall_211,ceiling_18]=True
    close[wall_211,shower_36]=True
    close[wall_211,toilet_37]=True
    close[wall_211,door_44]=True
    close[wall_211,doorjamb_45]=True
    close[wall_211,floor_77]=True
    close[wall_211,wall_84]=True
    close[wall_211,wall_85]=True
    close[wall_211,ceiling_95]=True
    close[wall_211,trashcan_99]=True
    close[wall_211,doorjamb_165]=True
    close[wall_211,drawing_174]=True
    close[wall_211,floor_202]=True
    close[wall_211,floor_203]=True
    close[wall_211,floor_204]=True
    close[wall_211,floor_206]=True
    close[wall_211,wall_209]=True
    close[wall_211,wall_212]=True
    close[wall_211,ceiling_216]=True
    close[wall_211,ceiling_217]=True
    close[wall_211,ceiling_221]=True
    close[wall_211,door_222]=True
    close[wall_211,ceilinglamp_224]=True
    close[wall_211,table_226]=True
    close[wall_211,bench_228]=True
    close[wall_211,cupboard_229]=True
    close[wall_211,kitchen_counter_230]=True
    close[wall_211,sink_231]=True
    close[wall_211,faucet_232]=True
    close[wall_211,mat_236]=True
    close[wall_211,mat_237]=True
    close[wall_211,drawing_238]=True
    close[wall_211,drawing_239]=True
    close[wall_211,drawing_240]=True
    close[wall_211,light_245]=True
    close[wall_211,powersocket_246]=True
    close[wall_211,phone_247]=True
    close[wall_211,wall_clock_249]=True
    close[wall_211,fridge_289]=True
    close[wall_211,coffe_maker_290]=True
    close[wall_211,toaster_292]=True
    close[wall_211,microwave_297]=True
    close[wall_212,wall_15]=True
    close[wall_212,shower_36]=True
    close[wall_212,toilet_37]=True
    close[wall_212,floor_202]=True
    close[wall_212,floor_203]=True
    close[wall_212,floor_204]=True
    close[wall_212,floor_205]=True
    close[wall_212,wall_211]=True
    close[wall_212,wall_214]=True
    close[wall_212,wall_215]=True
    close[wall_212,ceiling_216]=True
    close[wall_212,ceiling_220]=True
    close[wall_212,ceiling_221]=True
    close[wall_212,ceilinglamp_224]=True
    close[wall_212,table_226]=True
    close[wall_212,bench_228]=True
    close[wall_212,cupboard_229]=True
    close[wall_212,kitchen_counter_230]=True
    close[wall_212,sink_231]=True
    close[wall_212,faucet_232]=True
    close[wall_212,wallshelf_234]=True
    close[wall_212,mat_236]=True
    close[wall_212,mat_237]=True
    close[wall_212,drawing_241]=True
    close[wall_212,drawing_242]=True
    close[wall_212,drawing_243]=True
    close[wall_212,stovefan_288]=True
    close[wall_212,coffe_maker_290]=True
    close[wall_212,toaster_292]=True
    close[wall_212,oven_295]=True
    close[wall_212,tray_296]=True
    close[wall_212,microwave_297]=True
    close[wall_212,drawing_403]=True
    close[wall_212,photoframe_430]=True
    close[wall_213,floor_205]=True
    close[wall_213,floor_207]=True
    close[wall_213,floor_208]=True
    close[wall_213,wall_210]=True
    close[wall_213,wall_214]=True
    close[wall_213,ceiling_218]=True
    close[wall_213,ceiling_219]=True
    close[wall_213,ceiling_220]=True
    close[wall_213,ceilinglamp_223]=True
    close[wall_213,tvstand_225]=True
    close[wall_213,table_226]=True
    close[wall_213,bench_227]=True
    close[wall_213,wallshelf_235]=True
    close[wall_213,mat_236]=True
    close[wall_213,mat_237]=True
    close[wall_213,drawing_242]=True
    close[wall_213,orchid_244]=True
    close[wall_213,television_248]=True
    close[wall_213,photoframe_285]=True
    close[wall_213,floor_325]=True
    close[wall_213,wall_331]=True
    close[wall_213,ceiling_342]=True
    close[wall_213,doorjamb_346]=True
    close[wall_213,desk_357]=True
    close[wall_213,filing_cabinet_399]=True
    close[wall_213,drawing_402]=True
    close[wall_213,drawing_403]=True
    close[wall_213,drawing_404]=True
    close[wall_213,light_411]=True
    close[wall_213,powersocket_412]=True
    close[wall_213,mouse_413]=True
    close[wall_213,mousepad_414]=True
    close[wall_213,keyboard_415]=True
    close[wall_213,cpuscreen_416]=True
    close[wall_213,computer_417]=True
    close[wall_214,floor_205]=True
    close[wall_214,wall_212]=True
    close[wall_214,wall_213]=True
    close[wall_214,wall_215]=True
    close[wall_214,ceiling_220]=True
    close[wall_214,table_226]=True
    close[wall_214,wallshelf_234]=True
    close[wall_214,wallshelf_235]=True
    close[wall_214,mat_236]=True
    close[wall_214,drawing_241]=True
    close[wall_214,drawing_242]=True
    close[wall_214,drawing_243]=True
    close[wall_214,floor_320]=True
    close[wall_214,wall_331]=True
    close[wall_214,wall_332]=True
    close[wall_214,ceiling_337]=True
    close[wall_214,doorjamb_346]=True
    close[wall_214,bookshelf_354]=True
    close[wall_214,filing_cabinet_399]=True
    close[wall_214,drawing_402]=True
    close[wall_214,drawing_403]=True
    close[wall_214,drawing_404]=True
    close[wall_214,light_411]=True
    close[wall_214,photoframe_430]=True
    close[wall_215,floor_204]=True
    close[wall_215,wall_212]=True
    close[wall_215,wall_214]=True
    close[wall_215,ceiling_221]=True
    close[wall_215,wallshelf_234]=True
    close[wall_215,drawing_241]=True
    close[wall_215,drawing_242]=True
    close[wall_215,drawing_243]=True
    close[wall_215,stovefan_288]=True
    close[wall_215,coffe_maker_290]=True
    close[wall_215,oven_295]=True
    close[wall_215,tray_296]=True
    close[wall_215,floor_320]=True
    close[wall_215,wall_332]=True
    close[wall_215,wall_335]=True
    close[wall_215,ceiling_337]=True
    close[wall_215,walllamp_350]=True
    close[wall_215,bookshelf_354]=True
    close[wall_215,drawing_403]=True
    close[wall_215,photoframe_430]=True
    close[ceiling_216,wall_11]=True
    close[ceiling_216,ceiling_18]=True
    close[ceiling_216,shower_36]=True
    close[ceiling_216,wall_85]=True
    close[ceiling_216,ceiling_95]=True
    close[ceiling_216,drawing_174]=True
    close[ceiling_216,wall_211]=True
    close[ceiling_216,wall_212]=True
    close[ceiling_216,ceiling_217]=True
    close[ceiling_216,ceiling_221]=True
    close[ceiling_216,ceilinglamp_224]=True
    close[ceiling_216,cupboard_229]=True
    close[ceiling_216,faucet_232]=True
    close[ceiling_216,drawing_238]=True
    close[ceiling_216,drawing_239]=True
    close[ceiling_216,drawing_240]=True
    close[ceiling_216,light_245]=True
    close[ceiling_216,phone_247]=True
    close[ceiling_216,wall_clock_249]=True
    close[ceiling_216,fridge_289]=True
    close[ceiling_216,toaster_292]=True
    close[ceiling_216,microwave_297]=True
    close[ceiling_217,wall_84]=True
    close[ceiling_217,ceiling_94]=True
    close[ceiling_217,doorjamb_165]=True
    close[ceiling_217,light_169]=True
    close[ceiling_217,drawing_174]=True
    close[ceiling_217,wall_209]=True
    close[ceiling_217,wall_210]=True
    close[ceiling_217,wall_211]=True
    close[ceiling_217,ceiling_216]=True
    close[ceiling_217,ceiling_218]=True
    close[ceiling_217,ceiling_220]=True
    close[ceiling_217,ceilinglamp_223]=True
    close[ceiling_217,ceilinglamp_224]=True
    close[ceiling_217,drawing_238]=True
    close[ceiling_217,drawing_239]=True
    close[ceiling_217,drawing_240]=True
    close[ceiling_217,light_245]=True
    close[ceiling_217,phone_247]=True
    close[ceiling_217,wall_clock_249]=True
    close[ceiling_218,wall_83]=True
    close[ceiling_218,ceiling_93]=True
    close[ceiling_218,light_169]=True
    close[ceiling_218,cpuscreen_171]=True
    close[ceiling_218,wall_210]=True
    close[ceiling_218,wall_213]=True
    close[ceiling_218,ceiling_217]=True
    close[ceiling_218,ceiling_219]=True
    close[ceiling_218,ceilinglamp_223]=True
    close[ceiling_218,bookshelf_233]=True
    close[ceiling_219,wall_210]=True
    close[ceiling_219,wall_213]=True
    close[ceiling_219,ceiling_218]=True
    close[ceiling_219,ceiling_220]=True
    close[ceiling_219,ceilinglamp_223]=True
    close[ceiling_219,wallshelf_235]=True
    close[ceiling_219,wall_331]=True
    close[ceiling_219,ceiling_342]=True
    close[ceiling_219,doorjamb_346]=True
    close[ceiling_219,drawing_402]=True
    close[ceiling_219,drawing_404]=True
    close[ceiling_219,light_411]=True
    close[ceiling_220,wall_212]=True
    close[ceiling_220,wall_213]=True
    close[ceiling_220,wall_214]=True
    close[ceiling_220,ceiling_217]=True
    close[ceiling_220,ceiling_219]=True
    close[ceiling_220,ceiling_221]=True
    close[ceiling_220,ceilinglamp_223]=True
    close[ceiling_220,ceilinglamp_224]=True
    close[ceiling_220,wallshelf_234]=True
    close[ceiling_220,wallshelf_235]=True
    close[ceiling_220,drawing_241]=True
    close[ceiling_220,drawing_242]=True
    close[ceiling_220,drawing_243]=True
    close[ceiling_220,wall_332]=True
    close[ceiling_220,ceiling_337]=True
    close[ceiling_220,drawing_402]=True
    close[ceiling_220,drawing_403]=True
    close[ceiling_220,drawing_404]=True
    close[ceiling_220,light_411]=True
    close[ceiling_221,wall_15]=True
    close[ceiling_221,wall_211]=True
    close[ceiling_221,wall_212]=True
    close[ceiling_221,wall_215]=True
    close[ceiling_221,ceiling_216]=True
    close[ceiling_221,ceiling_220]=True
    close[ceiling_221,ceilinglamp_224]=True
    close[ceiling_221,cupboard_229]=True
    close[ceiling_221,faucet_232]=True
    close[ceiling_221,wallshelf_234]=True
    close[ceiling_221,drawing_241]=True
    close[ceiling_221,drawing_243]=True
    close[ceiling_221,stovefan_288]=True
    close[ceiling_221,coffe_maker_290]=True
    close[ceiling_221,toaster_292]=True
    close[ceiling_221,oven_295]=True
    close[ceiling_221,drawing_403]=True
    close[door_222,floor_75]=True
    close[door_222,floor_76]=True
    close[door_222,floor_77]=True
    close[door_222,wall_83]=True
    close[door_222,wall_84]=True
    close[door_222,wall_85]=True
    close[door_222,trashcan_99]=True
    close[door_222,desk_104]=True
    close[door_222,doorjamb_165]=True
    close[door_222,light_169]=True
    close[door_222,computer_170]=True
    close[door_222,drawing_174]=True
    close[door_222,floor_202]=True
    close[door_222,floor_203]=True
    close[door_222,floor_206]=True
    close[door_222,floor_207]=True
    close[door_222,wall_209]=True
    close[door_222,wall_210]=True
    close[door_222,wall_211]=True
    close[door_222,bookshelf_233]=True
    close[door_222,drawing_238]=True
    close[door_222,drawing_240]=True
    close[door_222,light_245]=True
    close[door_222,powersocket_246]=True
    close[door_222,phone_247]=True
    close[door_222,wall_clock_249]=True
    close[ceilinglamp_223,wall_210]=True
    close[ceilinglamp_223,wall_213]=True
    close[ceilinglamp_223,ceiling_217]=True
    close[ceilinglamp_223,ceiling_218]=True
    close[ceilinglamp_223,ceiling_219]=True
    close[ceilinglamp_223,ceiling_220]=True
    close[ceilinglamp_224,wall_211]=True
    close[ceilinglamp_224,wall_212]=True
    close[ceilinglamp_224,ceiling_216]=True
    close[ceilinglamp_224,ceiling_217]=True
    close[ceilinglamp_224,ceiling_220]=True
    close[ceilinglamp_224,ceiling_221]=True
    close[ceilinglamp_224,table_226]=True
    close[tvstand_225,cd_player_2060]=True
    close[tvstand_225,cd_2075]=True
    close[tvstand_225,floor_207]=True
    close[tvstand_225,floor_208]=True
    close[tvstand_225,wall_210]=True
    close[tvstand_225,wall_213]=True
    close[tvstand_225,orchid_244]=True
    close[tvstand_225,television_248]=True
    close[tvstand_225,photoframe_285]=True
    close[tvstand_225,powersocket_412]=True
    close[table_226,bowl_2071]=True
    close[table_226,bowl_2072]=True
    close[table_226,fork_2080]=True
    close[table_226,fork_2081]=True
    close[table_226,floor_202]=True
    close[table_226,floor_203]=True
    close[table_226,floor_204]=True
    close[table_226,floor_205]=True
    close[table_226,floor_206]=True
    close[table_226,floor_207]=True
    close[table_226,floor_208]=True
    close[table_226,wall_210]=True
    close[table_226,wall_211]=True
    close[table_226,wall_212]=True
    close[table_226,wall_213]=True
    close[table_226,wall_214]=True
    close[table_226,ceilinglamp_224]=True
    close[table_226,bench_227]=True
    close[table_226,bench_228]=True
    close[table_226,wallshelf_235]=True
    close[table_226,mat_236]=True
    close[table_226,mat_237]=True
    close[table_226,drawing_241]=True
    close[table_226,drawing_242]=True
    close[table_226,drawing_243]=True
    close[table_226,drawing_402]=True
    close[table_226,drawing_403]=True
    close[table_226,coffee_filter_2000]=True
    close[table_226,drawing_2003]=True
    close[bench_227,floor_205]=True
    close[bench_227,floor_206]=True
    close[bench_227,floor_207]=True
    close[bench_227,floor_208]=True
    close[bench_227,wall_210]=True
    close[bench_227,wall_213]=True
    close[bench_227,table_226]=True
    close[bench_227,bench_228]=True
    close[bench_227,mat_236]=True
    close[bench_227,mat_237]=True
    close[bench_228,floor_202]=True
    close[bench_228,floor_203]=True
    close[bench_228,floor_204]=True
    close[bench_228,floor_205]=True
    close[bench_228,floor_206]=True
    close[bench_228,wall_211]=True
    close[bench_228,wall_212]=True
    close[bench_228,table_226]=True
    close[bench_228,bench_227]=True
    close[bench_228,mat_236]=True
    close[bench_228,mat_237]=True
    close[cupboard_229,wall_11]=True
    close[cupboard_229,wall_15]=True
    close[cupboard_229,ceiling_18]=True
    close[cupboard_229,shower_36]=True
    close[cupboard_229,wall_211]=True
    close[cupboard_229,wall_212]=True
    close[cupboard_229,ceiling_216]=True
    close[cupboard_229,ceiling_221]=True
    close[cupboard_229,kitchen_counter_230]=True
    close[cupboard_229,sink_231]=True
    close[cupboard_229,faucet_232]=True
    close[cupboard_229,stovefan_288]=True
    close[cupboard_229,fridge_289]=True
    close[cupboard_229,coffe_maker_290]=True
    close[cupboard_229,toaster_292]=True
    close[cupboard_229,oven_295]=True
    close[cupboard_229,tray_296]=True
    close[cupboard_229,microwave_297]=True
    close[kitchen_counter_230,knife_2050]=True
    close[kitchen_counter_230,cutting_board_2051]=True
    close[kitchen_counter_230,cup_2063]=True
    close[kitchen_counter_230,cup_2064]=True
    close[kitchen_counter_230,stove_2065]=True
    close[kitchen_counter_230,pot_2069]=True
    close[kitchen_counter_230,oil_2079]=True
    close[kitchen_counter_230,fryingpan_2083]=True
    close[kitchen_counter_230,floor_7]=True
    close[kitchen_counter_230,wall_11]=True
    close[kitchen_counter_230,wall_15]=True
    close[kitchen_counter_230,shower_36]=True
    close[kitchen_counter_230,toilet_37]=True
    close[kitchen_counter_230,trashcan_99]=True
    close[kitchen_counter_230,drawing_174]=True
    close[kitchen_counter_230,floor_202]=True
    close[kitchen_counter_230,floor_203]=True
    close[kitchen_counter_230,floor_204]=True
    close[kitchen_counter_230,wall_211]=True
    close[kitchen_counter_230,wall_212]=True
    close[kitchen_counter_230,cupboard_229]=True
    close[kitchen_counter_230,sink_231]=True
    close[kitchen_counter_230,faucet_232]=True
    close[kitchen_counter_230,drawing_239]=True
    close[kitchen_counter_230,stovefan_288]=True
    close[kitchen_counter_230,fridge_289]=True
    close[kitchen_counter_230,coffe_maker_290]=True
    close[kitchen_counter_230,toaster_292]=True
    close[kitchen_counter_230,oven_295]=True
    close[kitchen_counter_230,tray_296]=True
    close[kitchen_counter_230,microwave_297]=True
    close[kitchen_counter_230,napkin_2005]=True
    close[sink_231,soap_2054]=True
    close[sink_231,floor_7]=True
    close[sink_231,wall_11]=True
    close[sink_231,wall_15]=True
    close[sink_231,shower_36]=True
    close[sink_231,toilet_37]=True
    close[sink_231,floor_202]=True
    close[sink_231,floor_203]=True
    close[sink_231,floor_204]=True
    close[sink_231,wall_211]=True
    close[sink_231,wall_212]=True
    close[sink_231,cupboard_229]=True
    close[sink_231,kitchen_counter_230]=True
    close[sink_231,faucet_232]=True
    close[sink_231,coffe_maker_290]=True
    close[sink_231,toaster_292]=True
    close[sink_231,microwave_297]=True
    close[sink_231,plate_1000]=True
    close[sink_231,dishwasher_1001]=True
    close[faucet_232,floor_7]=True
    close[faucet_232,wall_11]=True
    close[faucet_232,wall_15]=True
    close[faucet_232,ceiling_18]=True
    close[faucet_232,shower_36]=True
    close[faucet_232,toilet_37]=True
    close[faucet_232,floor_202]=True
    close[faucet_232,floor_203]=True
    close[faucet_232,floor_204]=True
    close[faucet_232,wall_211]=True
    close[faucet_232,wall_212]=True
    close[faucet_232,ceiling_216]=True
    close[faucet_232,ceiling_221]=True
    close[faucet_232,cupboard_229]=True
    close[faucet_232,kitchen_counter_230]=True
    close[faucet_232,sink_231]=True
    close[faucet_232,coffe_maker_290]=True
    close[faucet_232,toaster_292]=True
    close[faucet_232,oven_295]=True
    close[faucet_232,microwave_297]=True
    close[bookshelf_233,floor_75]=True
    close[bookshelf_233,floor_76]=True
    close[bookshelf_233,wall_83]=True
    close[bookshelf_233,wall_84]=True
    close[bookshelf_233,ceiling_93]=True
    close[bookshelf_233,chair_103]=True
    close[bookshelf_233,desk_104]=True
    close[bookshelf_233,doorjamb_165]=True
    close[bookshelf_233,mouse_166]=True
    close[bookshelf_233,mousepad_167]=True
    close[bookshelf_233,keyboard_168]=True
    close[bookshelf_233,light_169]=True
    close[bookshelf_233,computer_170]=True
    close[bookshelf_233,cpuscreen_171]=True
    close[bookshelf_233,floor_206]=True
    close[bookshelf_233,floor_207]=True
    close[bookshelf_233,wall_209]=True
    close[bookshelf_233,wall_210]=True
    close[bookshelf_233,ceiling_218]=True
    close[bookshelf_233,door_222]=True
    close[wallshelf_234,wall_212]=True
    close[wallshelf_234,wall_214]=True
    close[wallshelf_234,wall_215]=True
    close[wallshelf_234,ceiling_220]=True
    close[wallshelf_234,ceiling_221]=True
    close[wallshelf_234,drawing_241]=True
    close[wallshelf_234,drawing_242]=True
    close[wallshelf_234,drawing_243]=True
    close[wallshelf_234,stovefan_288]=True
    close[wallshelf_234,oven_295]=True
    close[wallshelf_234,wall_332]=True
    close[wallshelf_234,ceiling_337]=True
    close[wallshelf_234,bookshelf_354]=True
    close[wallshelf_234,drawing_403]=True
    close[wallshelf_234,photoframe_430]=True
    close[wallshelf_235,wall_213]=True
    close[wallshelf_235,wall_214]=True
    close[wallshelf_235,ceiling_219]=True
    close[wallshelf_235,ceiling_220]=True
    close[wallshelf_235,table_226]=True
    close[wallshelf_235,drawing_241]=True
    close[wallshelf_235,drawing_242]=True
    close[wallshelf_235,drawing_243]=True
    close[wallshelf_235,wall_331]=True
    close[wallshelf_235,wall_332]=True
    close[wallshelf_235,ceiling_337]=True
    close[wallshelf_235,ceiling_342]=True
    close[wallshelf_235,doorjamb_346]=True
    close[wallshelf_235,filing_cabinet_399]=True
    close[wallshelf_235,drawing_402]=True
    close[wallshelf_235,drawing_403]=True
    close[wallshelf_235,drawing_404]=True
    close[wallshelf_235,light_411]=True
    close[mat_236,floor_205]=True
    close[mat_236,floor_206]=True
    close[mat_236,wall_210]=True
    close[mat_236,wall_211]=True
    close[mat_236,wall_212]=True
    close[mat_236,wall_213]=True
    close[mat_236,wall_214]=True
    close[mat_236,table_226]=True
    close[mat_236,bench_227]=True
    close[mat_236,bench_228]=True
    close[mat_236,mat_237]=True
    close[mat_236,drawing_241]=True
    close[mat_236,drawing_242]=True
    close[mat_236,drawing_243]=True
    close[mat_237,floor_202]=True
    close[mat_237,floor_203]=True
    close[mat_237,floor_204]=True
    close[mat_237,floor_205]=True
    close[mat_237,floor_206]=True
    close[mat_237,floor_207]=True
    close[mat_237,floor_208]=True
    close[mat_237,wall_210]=True
    close[mat_237,wall_211]=True
    close[mat_237,wall_212]=True
    close[mat_237,wall_213]=True
    close[mat_237,table_226]=True
    close[mat_237,bench_227]=True
    close[mat_237,bench_228]=True
    close[mat_237,mat_236]=True
    close[mat_237,orchid_244]=True
    close[drawing_238,floor_76]=True
    close[drawing_238,floor_77]=True
    close[drawing_238,wall_84]=True
    close[drawing_238,wall_85]=True
    close[drawing_238,ceiling_94]=True
    close[drawing_238,ceiling_95]=True
    close[drawing_238,trashcan_99]=True
    close[drawing_238,doorjamb_165]=True
    close[drawing_238,drawing_174]=True
    close[drawing_238,floor_202]=True
    close[drawing_238,floor_203]=True
    close[drawing_238,floor_206]=True
    close[drawing_238,wall_209]=True
    close[drawing_238,wall_211]=True
    close[drawing_238,ceiling_216]=True
    close[drawing_238,ceiling_217]=True
    close[drawing_238,door_222]=True
    close[drawing_238,drawing_239]=True
    close[drawing_238,drawing_240]=True
    close[drawing_238,light_245]=True
    close[drawing_238,powersocket_246]=True
    close[drawing_238,phone_247]=True
    close[drawing_238,wall_clock_249]=True
    close[drawing_239,wall_84]=True
    close[drawing_239,wall_85]=True
    close[drawing_239,ceiling_94]=True
    close[drawing_239,ceiling_95]=True
    close[drawing_239,trashcan_99]=True
    close[drawing_239,drawing_174]=True
    close[drawing_239,floor_202]=True
    close[drawing_239,floor_203]=True
    close[drawing_239,wall_209]=True
    close[drawing_239,wall_211]=True
    close[drawing_239,ceiling_216]=True
    close[drawing_239,ceiling_217]=True
    close[drawing_239,kitchen_counter_230]=True
    close[drawing_239,drawing_238]=True
    close[drawing_239,drawing_240]=True
    close[drawing_239,light_245]=True
    close[drawing_239,phone_247]=True
    close[drawing_239,wall_clock_249]=True
    close[drawing_239,fridge_289]=True
    close[drawing_239,microwave_297]=True
    close[drawing_240,wall_84]=True
    close[drawing_240,wall_85]=True
    close[drawing_240,ceiling_94]=True
    close[drawing_240,ceiling_95]=True
    close[drawing_240,trashcan_99]=True
    close[drawing_240,doorjamb_165]=True
    close[drawing_240,drawing_174]=True
    close[drawing_240,wall_209]=True
    close[drawing_240,wall_211]=True
    close[drawing_240,ceiling_216]=True
    close[drawing_240,ceiling_217]=True
    close[drawing_240,door_222]=True
    close[drawing_240,drawing_238]=True
    close[drawing_240,drawing_239]=True
    close[drawing_240,light_245]=True
    close[drawing_240,phone_247]=True
    close[drawing_240,wall_clock_249]=True
    close[drawing_240,fridge_289]=True
    close[drawing_241,wall_212]=True
    close[drawing_241,wall_214]=True
    close[drawing_241,wall_215]=True
    close[drawing_241,ceiling_220]=True
    close[drawing_241,ceiling_221]=True
    close[drawing_241,table_226]=True
    close[drawing_241,wallshelf_234]=True
    close[drawing_241,wallshelf_235]=True
    close[drawing_241,mat_236]=True
    close[drawing_241,drawing_242]=True
    close[drawing_241,drawing_243]=True
    close[drawing_241,wall_332]=True
    close[drawing_241,ceiling_337]=True
    close[drawing_241,bookshelf_354]=True
    close[drawing_241,filing_cabinet_399]=True
    close[drawing_241,drawing_402]=True
    close[drawing_241,drawing_403]=True
    close[drawing_241,drawing_404]=True
    close[drawing_241,photoframe_430]=True
    close[drawing_242,floor_205]=True
    close[drawing_242,wall_212]=True
    close[drawing_242,wall_213]=True
    close[drawing_242,wall_214]=True
    close[drawing_242,wall_215]=True
    close[drawing_242,ceiling_220]=True
    close[drawing_242,table_226]=True
    close[drawing_242,wallshelf_234]=True
    close[drawing_242,wallshelf_235]=True
    close[drawing_242,mat_236]=True
    close[drawing_242,drawing_241]=True
    close[drawing_242,drawing_243]=True
    close[drawing_242,floor_320]=True
    close[drawing_242,wall_331]=True
    close[drawing_242,wall_332]=True
    close[drawing_242,ceiling_337]=True
    close[drawing_242,bookshelf_354]=True
    close[drawing_242,filing_cabinet_399]=True
    close[drawing_242,drawing_402]=True
    close[drawing_242,drawing_403]=True
    close[drawing_242,drawing_404]=True
    close[drawing_243,floor_204]=True
    close[drawing_243,floor_205]=True
    close[drawing_243,wall_212]=True
    close[drawing_243,wall_214]=True
    close[drawing_243,wall_215]=True
    close[drawing_243,ceiling_220]=True
    close[drawing_243,ceiling_221]=True
    close[drawing_243,table_226]=True
    close[drawing_243,wallshelf_234]=True
    close[drawing_243,wallshelf_235]=True
    close[drawing_243,mat_236]=True
    close[drawing_243,drawing_241]=True
    close[drawing_243,drawing_242]=True
    close[drawing_243,floor_320]=True
    close[drawing_243,wall_332]=True
    close[drawing_243,ceiling_337]=True
    close[drawing_243,bookshelf_354]=True
    close[drawing_243,filing_cabinet_399]=True
    close[drawing_243,drawing_402]=True
    close[drawing_243,drawing_403]=True
    close[drawing_243,drawing_404]=True
    close[drawing_243,photoframe_430]=True
    close[orchid_244,floor_207]=True
    close[orchid_244,floor_208]=True
    close[orchid_244,wall_210]=True
    close[orchid_244,wall_213]=True
    close[orchid_244,tvstand_225]=True
    close[orchid_244,mat_237]=True
    close[orchid_244,television_248]=True
    close[orchid_244,photoframe_285]=True
    close[light_245,floor_76]=True
    close[light_245,floor_77]=True
    close[light_245,wall_84]=True
    close[light_245,wall_85]=True
    close[light_245,ceiling_94]=True
    close[light_245,ceiling_95]=True
    close[light_245,trashcan_99]=True
    close[light_245,doorjamb_165]=True
    close[light_245,light_169]=True
    close[light_245,drawing_174]=True
    close[light_245,floor_202]=True
    close[light_245,floor_203]=True
    close[light_245,floor_206]=True
    close[light_245,wall_209]=True
    close[light_245,wall_211]=True
    close[light_245,ceiling_216]=True
    close[light_245,ceiling_217]=True
    close[light_245,door_222]=True
    close[light_245,drawing_238]=True
    close[light_245,drawing_239]=True
    close[light_245,drawing_240]=True
    close[light_245,powersocket_246]=True
    close[light_245,phone_247]=True
    close[light_245,wall_clock_249]=True
    close[powersocket_246,floor_76]=True
    close[powersocket_246,floor_77]=True
    close[powersocket_246,wall_84]=True
    close[powersocket_246,wall_85]=True
    close[powersocket_246,trashcan_99]=True
    close[powersocket_246,doorjamb_165]=True
    close[powersocket_246,light_169]=True
    close[powersocket_246,drawing_174]=True
    close[powersocket_246,floor_202]=True
    close[powersocket_246,floor_203]=True
    close[powersocket_246,floor_206]=True
    close[powersocket_246,wall_209]=True
    close[powersocket_246,wall_211]=True
    close[powersocket_246,door_222]=True
    close[powersocket_246,drawing_238]=True
    close[powersocket_246,light_245]=True
    close[powersocket_246,phone_247]=True
    close[phone_247,floor_76]=True
    close[phone_247,floor_77]=True
    close[phone_247,wall_84]=True
    close[phone_247,wall_85]=True
    close[phone_247,ceiling_94]=True
    close[phone_247,ceiling_95]=True
    close[phone_247,trashcan_99]=True
    close[phone_247,doorjamb_165]=True
    close[phone_247,light_169]=True
    close[phone_247,drawing_174]=True
    close[phone_247,floor_202]=True
    close[phone_247,floor_203]=True
    close[phone_247,floor_206]=True
    close[phone_247,wall_209]=True
    close[phone_247,wall_211]=True
    close[phone_247,ceiling_216]=True
    close[phone_247,ceiling_217]=True
    close[phone_247,door_222]=True
    close[phone_247,drawing_238]=True
    close[phone_247,drawing_239]=True
    close[phone_247,drawing_240]=True
    close[phone_247,light_245]=True
    close[phone_247,powersocket_246]=True
    close[phone_247,wall_clock_249]=True
    close[television_248,floor_207]=True
    close[television_248,floor_208]=True
    close[television_248,wall_210]=True
    close[television_248,wall_213]=True
    close[television_248,tvstand_225]=True
    close[television_248,orchid_244]=True
    close[television_248,photoframe_285]=True
    close[wall_clock_249,wall_84]=True
    close[wall_clock_249,wall_85]=True
    close[wall_clock_249,ceiling_94]=True
    close[wall_clock_249,ceiling_95]=True
    close[wall_clock_249,trashcan_99]=True
    close[wall_clock_249,doorjamb_165]=True
    close[wall_clock_249,drawing_174]=True
    close[wall_clock_249,wall_209]=True
    close[wall_clock_249,wall_211]=True
    close[wall_clock_249,ceiling_216]=True
    close[wall_clock_249,ceiling_217]=True
    close[wall_clock_249,door_222]=True
    close[wall_clock_249,drawing_238]=True
    close[wall_clock_249,drawing_239]=True
    close[wall_clock_249,drawing_240]=True
    close[wall_clock_249,light_245]=True
    close[wall_clock_249,phone_247]=True
    close[photoframe_285,floor_207]=True
    close[photoframe_285,floor_208]=True
    close[photoframe_285,wall_210]=True
    close[photoframe_285,wall_213]=True
    close[photoframe_285,tvstand_225]=True
    close[photoframe_285,orchid_244]=True
    close[photoframe_285,television_248]=True
    close[stovefan_288,wall_15]=True
    close[stovefan_288,wall_212]=True
    close[stovefan_288,wall_215]=True
    close[stovefan_288,ceiling_221]=True
    close[stovefan_288,cupboard_229]=True
    close[stovefan_288,kitchen_counter_230]=True
    close[stovefan_288,wallshelf_234]=True
    close[stovefan_288,coffe_maker_290]=True
    close[stovefan_288,toaster_292]=True
    close[stovefan_288,oven_295]=True
    close[stovefan_288,tray_296]=True
    close[fridge_289,food_steak_2008]=True
    close[fridge_289,food_apple_2009]=True
    close[fridge_289,food_bacon_2010]=True
    close[fridge_289,food_banana_2011]=True
    close[fridge_289,food_bread_2012]=True
    close[fridge_289,food_cake_2013]=True
    close[fridge_289,food_carrot_2014]=True
    close[fridge_289,food_cereal_2015]=True
    close[fridge_289,food_cheese_2016]=True
    close[fridge_289,food_chicken_2017]=True
    close[fridge_289,food_dessert_2018]=True
    close[fridge_289,food_donut_2019]=True
    close[fridge_289,food_egg_2020]=True
    close[fridge_289,food_fish_2021]=True
    close[fridge_289,food_food_2022]=True
    close[fridge_289,food_fruit_2023]=True
    close[fridge_289,food_hamburger_2024]=True
    close[fridge_289,food_ice_cream_2025]=True
    close[fridge_289,food_jam_2026]=True
    close[fridge_289,food_kiwi_2027]=True
    close[fridge_289,food_lemon_2028]=True
    close[fridge_289,food_noodles_2029]=True
    close[fridge_289,food_oatmeal_2030]=True
    close[fridge_289,food_orange_2031]=True
    close[fridge_289,food_onion_2032]=True
    close[fridge_289,food_peanut_butter_2033]=True
    close[fridge_289,food_pizza_2034]=True
    close[fridge_289,food_potato_2035]=True
    close[fridge_289,food_rice_2036]=True
    close[fridge_289,food_salt_2037]=True
    close[fridge_289,food_snack_2038]=True
    close[fridge_289,food_sugar_2039]=True
    close[fridge_289,food_turkey_2040]=True
    close[fridge_289,food_vegetable_2041]=True
    close[fridge_289,dry_pasta_2042]=True
    close[fridge_289,milk_2043]=True
    close[fridge_289,sauce_2078]=True
    close[fridge_289,floor_6]=True
    close[fridge_289,floor_7]=True
    close[fridge_289,wall_11]=True
    close[fridge_289,wall_14]=True
    close[fridge_289,ceiling_18]=True
    close[fridge_289,mat_22]=True
    close[fridge_289,shower_36]=True
    close[fridge_289,toilet_37]=True
    close[fridge_289,door_44]=True
    close[fridge_289,doorjamb_45]=True
    close[fridge_289,floor_77]=True
    close[fridge_289,wall_85]=True
    close[fridge_289,ceiling_95]=True
    close[fridge_289,trashcan_99]=True
    close[fridge_289,drawing_174]=True
    close[fridge_289,floor_202]=True
    close[fridge_289,floor_203]=True
    close[fridge_289,wall_211]=True
    close[fridge_289,ceiling_216]=True
    close[fridge_289,cupboard_229]=True
    close[fridge_289,kitchen_counter_230]=True
    close[fridge_289,drawing_239]=True
    close[fridge_289,drawing_240]=True
    close[fridge_289,microwave_297]=True
    close[coffe_maker_290,wall_11]=True
    close[coffe_maker_290,wall_15]=True
    close[coffe_maker_290,shower_36]=True
    close[coffe_maker_290,floor_204]=True
    close[coffe_maker_290,wall_211]=True
    close[coffe_maker_290,wall_212]=True
    close[coffe_maker_290,wall_215]=True
    close[coffe_maker_290,ceiling_221]=True
    close[coffe_maker_290,cupboard_229]=True
    close[coffe_maker_290,kitchen_counter_230]=True
    close[coffe_maker_290,sink_231]=True
    close[coffe_maker_290,faucet_232]=True
    close[coffe_maker_290,stovefan_288]=True
    close[coffe_maker_290,toaster_292]=True
    close[coffe_maker_290,oven_295]=True
    close[coffe_maker_290,tray_296]=True
    close[toaster_292,floor_7]=True
    close[toaster_292,wall_11]=True
    close[toaster_292,wall_15]=True
    close[toaster_292,shower_36]=True
    close[toaster_292,toilet_37]=True
    close[toaster_292,floor_202]=True
    close[toaster_292,floor_203]=True
    close[toaster_292,floor_204]=True
    close[toaster_292,wall_211]=True
    close[toaster_292,wall_212]=True
    close[toaster_292,ceiling_216]=True
    close[toaster_292,ceiling_221]=True
    close[toaster_292,cupboard_229]=True
    close[toaster_292,kitchen_counter_230]=True
    close[toaster_292,sink_231]=True
    close[toaster_292,faucet_232]=True
    close[toaster_292,stovefan_288]=True
    close[toaster_292,coffe_maker_290]=True
    close[toaster_292,oven_295]=True
    close[toaster_292,tray_296]=True
    close[toaster_292,microwave_297]=True
    close[oven_295,wall_15]=True
    close[oven_295,floor_204]=True
    close[oven_295,wall_212]=True
    close[oven_295,wall_215]=True
    close[oven_295,ceiling_221]=True
    close[oven_295,cupboard_229]=True
    close[oven_295,kitchen_counter_230]=True
    close[oven_295,faucet_232]=True
    close[oven_295,wallshelf_234]=True
    close[oven_295,stovefan_288]=True
    close[oven_295,coffe_maker_290]=True
    close[oven_295,toaster_292]=True
    close[oven_295,tray_296]=True
    close[tray_296,wall_15]=True
    close[tray_296,floor_204]=True
    close[tray_296,wall_212]=True
    close[tray_296,wall_215]=True
    close[tray_296,cupboard_229]=True
    close[tray_296,kitchen_counter_230]=True
    close[tray_296,stovefan_288]=True
    close[tray_296,coffe_maker_290]=True
    close[tray_296,toaster_292]=True
    close[tray_296,oven_295]=True
    close[microwave_297,floor_7]=True
    close[microwave_297,wall_11]=True
    close[microwave_297,wall_14]=True
    close[microwave_297,wall_15]=True
    close[microwave_297,ceiling_18]=True
    close[microwave_297,shower_36]=True
    close[microwave_297,toilet_37]=True
    close[microwave_297,wall_85]=True
    close[microwave_297,drawing_174]=True
    close[microwave_297,floor_202]=True
    close[microwave_297,floor_203]=True
    close[microwave_297,wall_211]=True
    close[microwave_297,wall_212]=True
    close[microwave_297,ceiling_216]=True
    close[microwave_297,cupboard_229]=True
    close[microwave_297,kitchen_counter_230]=True
    close[microwave_297,sink_231]=True
    close[microwave_297,faucet_232]=True
    close[microwave_297,drawing_239]=True
    close[microwave_297,fridge_289]=True
    close[microwave_297,toaster_292]=True
    close[home_office_319,coffee_table_2068]=True
    close[floor_320,floor_205]=True
    close[floor_320,wall_214]=True
    close[floor_320,wall_215]=True
    close[floor_320,drawing_242]=True
    close[floor_320,drawing_243]=True
    close[floor_320,floor_321]=True
    close[floor_320,floor_325]=True
    close[floor_320,wall_332]=True
    close[floor_320,bookshelf_354]=True
    close[floor_320,filing_cabinet_399]=True
    close[floor_320,light_411]=True
    close[floor_320,photoframe_430]=True
    close[floor_321,floor_320]=True
    close[floor_321,floor_322]=True
    close[floor_321,floor_324]=True
    close[floor_321,wall_332]=True
    close[floor_321,wall_333]=True
    close[floor_321,wall_335]=True
    close[floor_321,walllamp_350]=True
    close[floor_321,couch_352]=True
    close[floor_321,bookshelf_354]=True
    close[floor_321,table_355]=True
    close[floor_321,mat_401]=True
    close[floor_321,pillow_406]=True
    close[floor_322,floor_321]=True
    close[floor_322,floor_323]=True
    close[floor_322,wall_333]=True
    close[floor_322,couch_352]=True
    close[floor_322,table_355]=True
    close[floor_322,mat_401]=True
    close[floor_322,pillow_405]=True
    close[floor_322,pillow_406]=True
    close[floor_323,floor_322]=True
    close[floor_323,floor_324]=True
    close[floor_323,floor_328]=True
    close[floor_323,wall_329]=True
    close[floor_323,wall_333]=True
    close[floor_323,wall_334]=True
    close[floor_323,window_348]=True
    close[floor_323,couch_352]=True
    close[floor_323,tvstand_353]=True
    close[floor_323,table_355]=True
    close[floor_323,mat_401]=True
    close[floor_323,pillow_405]=True
    close[floor_323,curtain_407]=True
    close[floor_323,curtain_408]=True
    close[floor_323,curtain_409]=True
    close[floor_323,television_410]=True
    close[floor_324,floor_321]=True
    close[floor_324,floor_323]=True
    close[floor_324,floor_325]=True
    close[floor_324,floor_327]=True
    close[floor_324,couch_352]=True
    close[floor_324,tvstand_353]=True
    close[floor_324,table_355]=True
    close[floor_324,chair_356]=True
    close[floor_324,mat_401]=True
    close[floor_324,television_410]=True
    close[floor_325,floor_208]=True
    close[floor_325,wall_213]=True
    close[floor_325,floor_320]=True
    close[floor_325,floor_324]=True
    close[floor_325,floor_326]=True
    close[floor_325,wall_330]=True
    close[floor_325,wall_331]=True
    close[floor_325,wall_332]=True
    close[floor_325,doorjamb_346]=True
    close[floor_325,chair_356]=True
    close[floor_325,desk_357]=True
    close[floor_325,filing_cabinet_399]=True
    close[floor_325,light_411]=True
    close[floor_325,powersocket_412]=True
    close[floor_325,mouse_413]=True
    close[floor_325,mousepad_414]=True
    close[floor_325,keyboard_415]=True
    close[floor_325,computer_417]=True
    close[floor_326,floor_325]=True
    close[floor_326,floor_327]=True
    close[floor_326,wall_330]=True
    close[floor_326,walllamp_351]=True
    close[floor_326,chair_356]=True
    close[floor_326,desk_357]=True
    close[floor_326,powersocket_412]=True
    close[floor_326,mouse_413]=True
    close[floor_326,mousepad_414]=True
    close[floor_326,keyboard_415]=True
    close[floor_326,cpuscreen_416]=True
    close[floor_326,computer_417]=True
    close[floor_327,floor_324]=True
    close[floor_327,floor_326]=True
    close[floor_327,floor_328]=True
    close[floor_327,wall_330]=True
    close[floor_327,wall_334]=True
    close[floor_327,wall_336]=True
    close[floor_327,doorjamb_347]=True
    close[floor_327,walllamp_351]=True
    close[floor_327,tvstand_353]=True
    close[floor_327,chair_356]=True
    close[floor_327,dresser_358]=True
    close[floor_327,closetdrawer_377]=True
    close[floor_327,closetdrawer_380]=True
    close[floor_327,closetdrawer_382]=True
    close[floor_327,closetdrawer_384]=True
    close[floor_327,closetdrawer_388]=True
    close[floor_327,closetdrawer_392]=True
    close[floor_327,closetdrawer_394]=True
    close[floor_327,television_410]=True
    close[floor_328,floor_323]=True
    close[floor_328,floor_327]=True
    close[floor_328,wall_334]=True
    close[floor_328,tvstand_353]=True
    close[floor_328,dresser_358]=True
    close[floor_328,closetdrawer_377]=True
    close[floor_328,closetdrawer_380]=True
    close[floor_328,closetdrawer_382]=True
    close[floor_328,closetdrawer_384]=True
    close[floor_328,closetdrawer_388]=True
    close[floor_328,closetdrawer_392]=True
    close[floor_328,closetdrawer_394]=True
    close[floor_328,television_410]=True
    close[wall_329,floor_323]=True
    close[wall_329,wall_333]=True
    close[wall_329,wall_334]=True
    close[wall_329,ceiling_340]=True
    close[wall_329,window_348]=True
    close[wall_329,couch_352]=True
    close[wall_329,mat_401]=True
    close[wall_329,pillow_405]=True
    close[wall_329,curtain_407]=True
    close[wall_329,curtain_408]=True
    close[wall_329,curtain_409]=True
    close[wall_330,floor_325]=True
    close[wall_330,floor_326]=True
    close[wall_330,floor_327]=True
    close[wall_330,wall_331]=True
    close[wall_330,wall_336]=True
    close[wall_330,ceiling_342]=True
    close[wall_330,ceiling_343]=True
    close[wall_330,ceiling_344]=True
    close[wall_330,doorjamb_346]=True
    close[wall_330,doorjamb_347]=True
    close[wall_330,walllamp_351]=True
    close[wall_330,chair_356]=True
    close[wall_330,desk_357]=True
    close[wall_330,powersocket_412]=True
    close[wall_330,mouse_413]=True
    close[wall_330,mousepad_414]=True
    close[wall_330,keyboard_415]=True
    close[wall_330,cpuscreen_416]=True
    close[wall_330,computer_417]=True
    close[wall_331,floor_208]=True
    close[wall_331,wall_213]=True
    close[wall_331,wall_214]=True
    close[wall_331,ceiling_219]=True
    close[wall_331,wallshelf_235]=True
    close[wall_331,drawing_242]=True
    close[wall_331,floor_325]=True
    close[wall_331,wall_330]=True
    close[wall_331,wall_332]=True
    close[wall_331,ceiling_342]=True
    close[wall_331,doorjamb_346]=True
    close[wall_331,desk_357]=True
    close[wall_331,filing_cabinet_399]=True
    close[wall_331,drawing_402]=True
    close[wall_331,drawing_403]=True
    close[wall_331,drawing_404]=True
    close[wall_331,light_411]=True
    close[wall_331,powersocket_412]=True
    close[wall_331,mouse_413]=True
    close[wall_331,mousepad_414]=True
    close[wall_331,keyboard_415]=True
    close[wall_331,cpuscreen_416]=True
    close[wall_331,computer_417]=True
    close[wall_332,floor_205]=True
    close[wall_332,wall_214]=True
    close[wall_332,wall_215]=True
    close[wall_332,ceiling_220]=True
    close[wall_332,wallshelf_234]=True
    close[wall_332,wallshelf_235]=True
    close[wall_332,drawing_241]=True
    close[wall_332,drawing_242]=True
    close[wall_332,drawing_243]=True
    close[wall_332,floor_320]=True
    close[wall_332,floor_321]=True
    close[wall_332,floor_325]=True
    close[wall_332,wall_331]=True
    close[wall_332,wall_335]=True
    close[wall_332,ceiling_337]=True
    close[wall_332,ceiling_338]=True
    close[wall_332,ceiling_342]=True
    close[wall_332,doorjamb_346]=True
    close[wall_332,walllamp_350]=True
    close[wall_332,bookshelf_354]=True
    close[wall_332,filing_cabinet_399]=True
    close[wall_332,drawing_402]=True
    close[wall_332,drawing_403]=True
    close[wall_332,drawing_404]=True
    close[wall_332,light_411]=True
    close[wall_332,photoframe_430]=True
    close[wall_333,floor_321]=True
    close[wall_333,floor_322]=True
    close[wall_333,floor_323]=True
    close[wall_333,wall_329]=True
    close[wall_333,wall_335]=True
    close[wall_333,ceiling_338]=True
    close[wall_333,ceiling_339]=True
    close[wall_333,ceiling_340]=True
    close[wall_333,window_348]=True
    close[wall_333,couch_352]=True
    close[wall_333,table_355]=True
    close[wall_333,drawing_400]=True
    close[wall_333,mat_401]=True
    close[wall_333,pillow_405]=True
    close[wall_333,pillow_406]=True
    close[wall_333,curtain_409]=True
    close[wall_334,floor_323]=True
    close[wall_334,floor_327]=True
    close[wall_334,floor_328]=True
    close[wall_334,wall_329]=True
    close[wall_334,wall_336]=True
    close[wall_334,ceiling_340]=True
    close[wall_334,ceiling_344]=True
    close[wall_334,ceiling_345]=True
    close[wall_334,doorjamb_347]=True
    close[wall_334,window_348]=True
    close[wall_334,tvstand_353]=True
    close[wall_334,dresser_358]=True
    close[wall_334,hanger_359]=True
    close[wall_334,hanger_361]=True
    close[wall_334,hanger_363]=True
    close[wall_334,hanger_365]=True
    close[wall_334,hanger_367]=True
    close[wall_334,hanger_369]=True
    close[wall_334,hanger_372]=True
    close[wall_334,hanger_374]=True
    close[wall_334,hanger_375]=True
    close[wall_334,hanger_376]=True
    close[wall_334,closetdrawer_377]=True
    close[wall_334,closetdrawer_380]=True
    close[wall_334,closetdrawer_382]=True
    close[wall_334,closetdrawer_384]=True
    close[wall_334,closetdrawer_388]=True
    close[wall_334,closetdrawer_392]=True
    close[wall_334,closetdrawer_394]=True
    close[wall_334,curtain_407]=True
    close[wall_334,curtain_408]=True
    close[wall_334,television_410]=True
    close[wall_335,wall_215]=True
    close[wall_335,floor_321]=True
    close[wall_335,wall_332]=True
    close[wall_335,wall_333]=True
    close[wall_335,ceiling_338]=True
    close[wall_335,walllamp_350]=True
    close[wall_335,couch_352]=True
    close[wall_335,bookshelf_354]=True
    close[wall_335,drawing_400]=True
    close[wall_335,mat_401]=True
    close[wall_335,pillow_406]=True
    close[wall_335,photoframe_430]=True
    close[wall_336,floor_327]=True
    close[wall_336,wall_330]=True
    close[wall_336,wall_334]=True
    close[wall_336,ceiling_344]=True
    close[wall_336,doorjamb_347]=True
    close[wall_336,walllamp_351]=True
    close[wall_336,dresser_358]=True
    close[wall_336,hanger_359]=True
    close[wall_336,hanger_361]=True
    close[wall_336,hanger_363]=True
    close[wall_336,hanger_365]=True
    close[wall_336,hanger_367]=True
    close[wall_336,hanger_369]=True
    close[wall_336,hanger_372]=True
    close[wall_336,hanger_374]=True
    close[wall_336,hanger_375]=True
    close[wall_336,hanger_376]=True
    close[wall_336,closetdrawer_377]=True
    close[wall_336,closetdrawer_380]=True
    close[wall_336,closetdrawer_382]=True
    close[wall_336,closetdrawer_384]=True
    close[wall_336,closetdrawer_388]=True
    close[wall_336,closetdrawer_392]=True
    close[wall_336,closetdrawer_394]=True
    close[ceiling_337,wall_214]=True
    close[ceiling_337,wall_215]=True
    close[ceiling_337,ceiling_220]=True
    close[ceiling_337,wallshelf_234]=True
    close[ceiling_337,wallshelf_235]=True
    close[ceiling_337,drawing_241]=True
    close[ceiling_337,drawing_242]=True
    close[ceiling_337,drawing_243]=True
    close[ceiling_337,wall_332]=True
    close[ceiling_337,ceiling_338]=True
    close[ceiling_337,ceiling_342]=True
    close[ceiling_337,walllamp_350]=True
    close[ceiling_337,bookshelf_354]=True
    close[ceiling_337,drawing_402]=True
    close[ceiling_337,drawing_403]=True
    close[ceiling_337,drawing_404]=True
    close[ceiling_337,light_411]=True
    close[ceiling_337,photoframe_430]=True
    close[ceiling_338,wall_332]=True
    close[ceiling_338,wall_333]=True
    close[ceiling_338,wall_335]=True
    close[ceiling_338,ceiling_337]=True
    close[ceiling_338,ceiling_339]=True
    close[ceiling_338,ceiling_341]=True
    close[ceiling_338,ceilinglamp_349]=True
    close[ceiling_338,walllamp_350]=True
    close[ceiling_338,bookshelf_354]=True
    close[ceiling_338,drawing_400]=True
    close[ceiling_339,wall_333]=True
    close[ceiling_339,ceiling_338]=True
    close[ceiling_339,ceiling_340]=True
    close[ceiling_339,drawing_400]=True
    close[ceiling_339,curtain_409]=True
    close[ceiling_340,wall_329]=True
    close[ceiling_340,wall_333]=True
    close[ceiling_340,wall_334]=True
    close[ceiling_340,ceiling_339]=True
    close[ceiling_340,ceiling_341]=True
    close[ceiling_340,ceiling_345]=True
    close[ceiling_340,window_348]=True
    close[ceiling_340,ceilinglamp_349]=True
    close[ceiling_340,curtain_407]=True
    close[ceiling_340,curtain_408]=True
    close[ceiling_340,curtain_409]=True
    close[ceiling_340,television_410]=True
    close[ceiling_341,ceiling_338]=True
    close[ceiling_341,ceiling_340]=True
    close[ceiling_341,ceiling_342]=True
    close[ceiling_341,ceiling_344]=True
    close[ceiling_341,ceilinglamp_349]=True
    close[ceiling_341,television_410]=True
    close[ceiling_342,wall_213]=True
    close[ceiling_342,ceiling_219]=True
    close[ceiling_342,wallshelf_235]=True
    close[ceiling_342,wall_330]=True
    close[ceiling_342,wall_331]=True
    close[ceiling_342,wall_332]=True
    close[ceiling_342,ceiling_337]=True
    close[ceiling_342,ceiling_341]=True
    close[ceiling_342,ceiling_343]=True
    close[ceiling_342,doorjamb_346]=True
    close[ceiling_342,ceilinglamp_349]=True
    close[ceiling_342,drawing_402]=True
    close[ceiling_342,drawing_404]=True
    close[ceiling_342,light_411]=True
    close[ceiling_343,wall_330]=True
    close[ceiling_343,ceiling_342]=True
    close[ceiling_343,ceiling_344]=True
    close[ceiling_343,walllamp_351]=True
    close[ceiling_343,chair_356]=True
    close[ceiling_343,cpuscreen_416]=True
    close[ceiling_344,wall_330]=True
    close[ceiling_344,wall_334]=True
    close[ceiling_344,wall_336]=True
    close[ceiling_344,ceiling_341]=True
    close[ceiling_344,ceiling_343]=True
    close[ceiling_344,ceiling_345]=True
    close[ceiling_344,doorjamb_347]=True
    close[ceiling_344,ceilinglamp_349]=True
    close[ceiling_344,walllamp_351]=True
    close[ceiling_344,dresser_358]=True
    close[ceiling_344,hanger_359]=True
    close[ceiling_344,hanger_361]=True
    close[ceiling_344,hanger_363]=True
    close[ceiling_344,hanger_365]=True
    close[ceiling_344,hanger_369]=True
    close[ceiling_344,hanger_372]=True
    close[ceiling_344,hanger_374]=True
    close[ceiling_344,hanger_375]=True
    close[ceiling_344,hanger_376]=True
    close[ceiling_345,wall_334]=True
    close[ceiling_345,ceiling_340]=True
    close[ceiling_345,ceiling_344]=True
    close[ceiling_345,dresser_358]=True
    close[ceiling_345,hanger_359]=True
    close[ceiling_345,hanger_361]=True
    close[ceiling_345,hanger_363]=True
    close[ceiling_345,hanger_365]=True
    close[ceiling_345,hanger_367]=True
    close[ceiling_345,hanger_369]=True
    close[ceiling_345,hanger_372]=True
    close[ceiling_345,hanger_374]=True
    close[ceiling_345,hanger_375]=True
    close[ceiling_345,hanger_376]=True
    close[ceiling_345,curtain_407]=True
    close[ceiling_345,curtain_408]=True
    close[doorjamb_346,floor_208]=True
    close[doorjamb_346,wall_213]=True
    close[doorjamb_346,wall_214]=True
    close[doorjamb_346,ceiling_219]=True
    close[doorjamb_346,wallshelf_235]=True
    close[doorjamb_346,floor_325]=True
    close[doorjamb_346,wall_330]=True
    close[doorjamb_346,wall_331]=True
    close[doorjamb_346,wall_332]=True
    close[doorjamb_346,ceiling_342]=True
    close[doorjamb_346,desk_357]=True
    close[doorjamb_346,filing_cabinet_399]=True
    close[doorjamb_346,drawing_402]=True
    close[doorjamb_346,drawing_404]=True
    close[doorjamb_346,light_411]=True
    close[doorjamb_346,powersocket_412]=True
    close[doorjamb_346,mouse_413]=True
    close[doorjamb_346,mousepad_414]=True
    close[doorjamb_346,computer_417]=True
    close[doorjamb_347,floor_327]=True
    close[doorjamb_347,wall_330]=True
    close[doorjamb_347,wall_334]=True
    close[doorjamb_347,wall_336]=True
    close[doorjamb_347,ceiling_344]=True
    close[doorjamb_347,walllamp_351]=True
    close[doorjamb_347,dresser_358]=True
    close[doorjamb_347,hanger_359]=True
    close[doorjamb_347,hanger_374]=True
    close[doorjamb_347,hanger_375]=True
    close[doorjamb_347,hanger_376]=True
    close[doorjamb_347,closetdrawer_380]=True
    close[doorjamb_347,closetdrawer_382]=True
    close[doorjamb_347,closetdrawer_392]=True
    close[window_348,floor_323]=True
    close[window_348,wall_329]=True
    close[window_348,wall_333]=True
    close[window_348,wall_334]=True
    close[window_348,ceiling_340]=True
    close[window_348,couch_352]=True
    close[window_348,mat_401]=True
    close[window_348,pillow_405]=True
    close[window_348,curtain_407]=True
    close[window_348,curtain_408]=True
    close[window_348,curtain_409]=True
    close[ceilinglamp_349,ceiling_338]=True
    close[ceilinglamp_349,ceiling_340]=True
    close[ceilinglamp_349,ceiling_341]=True
    close[ceilinglamp_349,ceiling_342]=True
    close[ceilinglamp_349,ceiling_344]=True
    close[ceilinglamp_349,couch_352]=True
    close[ceilinglamp_349,television_410]=True
    close[walllamp_350,wall_215]=True
    close[walllamp_350,floor_321]=True
    close[walllamp_350,wall_332]=True
    close[walllamp_350,wall_335]=True
    close[walllamp_350,ceiling_337]=True
    close[walllamp_350,ceiling_338]=True
    close[walllamp_350,couch_352]=True
    close[walllamp_350,bookshelf_354]=True
    close[walllamp_350,mat_401]=True
    close[walllamp_350,pillow_406]=True
    close[walllamp_351,floor_326]=True
    close[walllamp_351,floor_327]=True
    close[walllamp_351,wall_330]=True
    close[walllamp_351,wall_336]=True
    close[walllamp_351,ceiling_343]=True
    close[walllamp_351,ceiling_344]=True
    close[walllamp_351,doorjamb_347]=True
    close[walllamp_351,chair_356]=True
    close[walllamp_351,desk_357]=True
    close[walllamp_351,keyboard_415]=True
    close[couch_352,clothes_jacket_2047]=True
    close[couch_352,remote_control_2052]=True
    close[couch_352,cat_2055]=True
    close[couch_352,vacuum_cleaner_2070]=True
    close[couch_352,floor_321]=True
    close[couch_352,floor_322]=True
    close[couch_352,floor_323]=True
    close[couch_352,floor_324]=True
    close[couch_352,wall_329]=True
    close[couch_352,wall_333]=True
    close[couch_352,wall_335]=True
    close[couch_352,window_348]=True
    close[couch_352,ceilinglamp_349]=True
    close[couch_352,walllamp_350]=True
    close[couch_352,tvstand_353]=True
    close[couch_352,table_355]=True
    close[couch_352,drawing_400]=True
    close[couch_352,mat_401]=True
    close[couch_352,pillow_405]=True
    close[couch_352,pillow_406]=True
    close[couch_352,curtain_407]=True
    close[couch_352,curtain_408]=True
    close[couch_352,curtain_409]=True
    close[couch_352,television_410]=True
    close[couch_352,hairbrush_2002]=True
    close[tvstand_353,dvd_player_2061]=True
    close[tvstand_353,floor_323]=True
    close[tvstand_353,floor_324]=True
    close[tvstand_353,floor_327]=True
    close[tvstand_353,floor_328]=True
    close[tvstand_353,wall_334]=True
    close[tvstand_353,couch_352]=True
    close[tvstand_353,table_355]=True
    close[tvstand_353,mat_401]=True
    close[tvstand_353,television_410]=True
    close[bookshelf_354,book_2066]=True
    close[bookshelf_354,book_2067]=True
    close[bookshelf_354,wall_214]=True
    close[bookshelf_354,wall_215]=True
    close[bookshelf_354,wallshelf_234]=True
    close[bookshelf_354,drawing_241]=True
    close[bookshelf_354,drawing_242]=True
    close[bookshelf_354,drawing_243]=True
    close[bookshelf_354,floor_320]=True
    close[bookshelf_354,floor_321]=True
    close[bookshelf_354,wall_332]=True
    close[bookshelf_354,wall_335]=True
    close[bookshelf_354,ceiling_337]=True
    close[bookshelf_354,ceiling_338]=True
    close[bookshelf_354,walllamp_350]=True
    close[bookshelf_354,filing_cabinet_399]=True
    close[bookshelf_354,drawing_402]=True
    close[bookshelf_354,drawing_403]=True
    close[bookshelf_354,photoframe_430]=True
    close[table_355,headset_2062]=True
    close[table_355,spectacles_2082]=True
    close[table_355,floor_321]=True
    close[table_355,floor_322]=True
    close[table_355,floor_323]=True
    close[table_355,floor_324]=True
    close[table_355,wall_333]=True
    close[table_355,couch_352]=True
    close[table_355,tvstand_353]=True
    close[table_355,mat_401]=True
    close[table_355,pillow_406]=True
    close[table_355,television_410]=True
    close[chair_356,floor_324]=True
    close[chair_356,floor_325]=True
    close[chair_356,floor_326]=True
    close[chair_356,floor_327]=True
    close[chair_356,wall_330]=True
    close[chair_356,ceiling_343]=True
    close[chair_356,walllamp_351]=True
    close[chair_356,desk_357]=True
    close[chair_356,mouse_413]=True
    close[chair_356,mousepad_414]=True
    close[chair_356,keyboard_415]=True
    close[chair_356,cpuscreen_416]=True
    close[chair_356,computer_417]=True
    close[desk_357,headset_2076]=True
    close[desk_357,phone_2077]=True
    close[desk_357,floor_208]=True
    close[desk_357,wall_213]=True
    close[desk_357,floor_325]=True
    close[desk_357,floor_326]=True
    close[desk_357,wall_330]=True
    close[desk_357,wall_331]=True
    close[desk_357,doorjamb_346]=True
    close[desk_357,walllamp_351]=True
    close[desk_357,chair_356]=True
    close[desk_357,powersocket_412]=True
    close[desk_357,mouse_413]=True
    close[desk_357,mousepad_414]=True
    close[desk_357,keyboard_415]=True
    close[desk_357,cpuscreen_416]=True
    close[desk_357,computer_417]=True
    close[desk_357,pencil_2001]=True
    close[dresser_358,floor_327]=True
    close[dresser_358,floor_328]=True
    close[dresser_358,wall_334]=True
    close[dresser_358,wall_336]=True
    close[dresser_358,ceiling_344]=True
    close[dresser_358,ceiling_345]=True
    close[dresser_358,doorjamb_347]=True
    close[dresser_358,hanger_359]=True
    close[dresser_358,hanger_361]=True
    close[dresser_358,hanger_363]=True
    close[dresser_358,hanger_365]=True
    close[dresser_358,hanger_367]=True
    close[dresser_358,hanger_369]=True
    close[dresser_358,hanger_372]=True
    close[dresser_358,hanger_374]=True
    close[dresser_358,hanger_375]=True
    close[dresser_358,hanger_376]=True
    close[dresser_358,closetdrawer_377]=True
    close[dresser_358,closetdrawer_380]=True
    close[dresser_358,closetdrawer_382]=True
    close[dresser_358,closetdrawer_384]=True
    close[dresser_358,closetdrawer_388]=True
    close[dresser_358,closetdrawer_392]=True
    close[dresser_358,closetdrawer_394]=True
    close[hanger_359,wall_334]=True
    close[hanger_359,wall_336]=True
    close[hanger_359,ceiling_344]=True
    close[hanger_359,ceiling_345]=True
    close[hanger_359,doorjamb_347]=True
    close[hanger_359,dresser_358]=True
    close[hanger_359,hanger_361]=True
    close[hanger_359,hanger_363]=True
    close[hanger_359,hanger_365]=True
    close[hanger_359,hanger_367]=True
    close[hanger_359,hanger_369]=True
    close[hanger_359,hanger_372]=True
    close[hanger_359,hanger_374]=True
    close[hanger_359,hanger_375]=True
    close[hanger_359,hanger_376]=True
    close[hanger_359,closetdrawer_377]=True
    close[hanger_359,closetdrawer_380]=True
    close[hanger_359,closetdrawer_382]=True
    close[hanger_359,closetdrawer_384]=True
    close[hanger_359,closetdrawer_388]=True
    close[hanger_361,wall_334]=True
    close[hanger_361,wall_336]=True
    close[hanger_361,ceiling_344]=True
    close[hanger_361,ceiling_345]=True
    close[hanger_361,dresser_358]=True
    close[hanger_361,hanger_359]=True
    close[hanger_361,hanger_363]=True
    close[hanger_361,hanger_365]=True
    close[hanger_361,hanger_367]=True
    close[hanger_361,hanger_369]=True
    close[hanger_361,hanger_372]=True
    close[hanger_361,hanger_374]=True
    close[hanger_361,hanger_375]=True
    close[hanger_361,hanger_376]=True
    close[hanger_361,closetdrawer_377]=True
    close[hanger_361,closetdrawer_380]=True
    close[hanger_361,closetdrawer_384]=True
    close[hanger_361,closetdrawer_388]=True
    close[hanger_363,wall_334]=True
    close[hanger_363,wall_336]=True
    close[hanger_363,ceiling_344]=True
    close[hanger_363,ceiling_345]=True
    close[hanger_363,dresser_358]=True
    close[hanger_363,hanger_359]=True
    close[hanger_363,hanger_361]=True
    close[hanger_363,hanger_365]=True
    close[hanger_363,hanger_367]=True
    close[hanger_363,hanger_369]=True
    close[hanger_363,hanger_372]=True
    close[hanger_363,hanger_374]=True
    close[hanger_363,hanger_375]=True
    close[hanger_363,hanger_376]=True
    close[hanger_363,closetdrawer_377]=True
    close[hanger_363,closetdrawer_380]=True
    close[hanger_363,closetdrawer_382]=True
    close[hanger_363,closetdrawer_384]=True
    close[hanger_363,closetdrawer_388]=True
    close[hanger_365,wall_334]=True
    close[hanger_365,wall_336]=True
    close[hanger_365,ceiling_344]=True
    close[hanger_365,ceiling_345]=True
    close[hanger_365,dresser_358]=True
    close[hanger_365,hanger_359]=True
    close[hanger_365,hanger_361]=True
    close[hanger_365,hanger_363]=True
    close[hanger_365,hanger_367]=True
    close[hanger_365,hanger_369]=True
    close[hanger_365,hanger_372]=True
    close[hanger_365,hanger_374]=True
    close[hanger_365,hanger_375]=True
    close[hanger_365,hanger_376]=True
    close[hanger_365,closetdrawer_377]=True
    close[hanger_365,closetdrawer_380]=True
    close[hanger_365,closetdrawer_382]=True
    close[hanger_365,closetdrawer_384]=True
    close[hanger_365,closetdrawer_388]=True
    close[hanger_367,wall_334]=True
    close[hanger_367,wall_336]=True
    close[hanger_367,ceiling_345]=True
    close[hanger_367,dresser_358]=True
    close[hanger_367,hanger_359]=True
    close[hanger_367,hanger_361]=True
    close[hanger_367,hanger_363]=True
    close[hanger_367,hanger_365]=True
    close[hanger_367,hanger_369]=True
    close[hanger_367,hanger_372]=True
    close[hanger_367,hanger_374]=True
    close[hanger_367,hanger_375]=True
    close[hanger_367,hanger_376]=True
    close[hanger_367,closetdrawer_377]=True
    close[hanger_367,closetdrawer_380]=True
    close[hanger_367,closetdrawer_384]=True
    close[hanger_367,closetdrawer_388]=True
    close[hanger_369,wall_334]=True
    close[hanger_369,wall_336]=True
    close[hanger_369,ceiling_344]=True
    close[hanger_369,ceiling_345]=True
    close[hanger_369,dresser_358]=True
    close[hanger_369,hanger_359]=True
    close[hanger_369,hanger_361]=True
    close[hanger_369,hanger_363]=True
    close[hanger_369,hanger_365]=True
    close[hanger_369,hanger_367]=True
    close[hanger_369,hanger_372]=True
    close[hanger_369,hanger_374]=True
    close[hanger_369,hanger_375]=True
    close[hanger_369,hanger_376]=True
    close[hanger_369,closetdrawer_377]=True
    close[hanger_369,closetdrawer_380]=True
    close[hanger_369,closetdrawer_384]=True
    close[hanger_369,closetdrawer_388]=True
    close[hanger_372,wall_334]=True
    close[hanger_372,wall_336]=True
    close[hanger_372,ceiling_344]=True
    close[hanger_372,ceiling_345]=True
    close[hanger_372,dresser_358]=True
    close[hanger_372,hanger_359]=True
    close[hanger_372,hanger_361]=True
    close[hanger_372,hanger_363]=True
    close[hanger_372,hanger_365]=True
    close[hanger_372,hanger_367]=True
    close[hanger_372,hanger_369]=True
    close[hanger_372,hanger_374]=True
    close[hanger_372,hanger_375]=True
    close[hanger_372,hanger_376]=True
    close[hanger_372,closetdrawer_377]=True
    close[hanger_372,closetdrawer_380]=True
    close[hanger_372,closetdrawer_382]=True
    close[hanger_372,closetdrawer_384]=True
    close[hanger_372,closetdrawer_388]=True
    close[hanger_374,wall_334]=True
    close[hanger_374,wall_336]=True
    close[hanger_374,ceiling_344]=True
    close[hanger_374,ceiling_345]=True
    close[hanger_374,doorjamb_347]=True
    close[hanger_374,dresser_358]=True
    close[hanger_374,hanger_359]=True
    close[hanger_374,hanger_361]=True
    close[hanger_374,hanger_363]=True
    close[hanger_374,hanger_365]=True
    close[hanger_374,hanger_367]=True
    close[hanger_374,hanger_369]=True
    close[hanger_374,hanger_372]=True
    close[hanger_374,hanger_375]=True
    close[hanger_374,hanger_376]=True
    close[hanger_374,closetdrawer_377]=True
    close[hanger_374,closetdrawer_380]=True
    close[hanger_374,closetdrawer_382]=True
    close[hanger_374,closetdrawer_384]=True
    close[hanger_374,closetdrawer_388]=True
    close[hanger_375,wall_334]=True
    close[hanger_375,wall_336]=True
    close[hanger_375,ceiling_344]=True
    close[hanger_375,ceiling_345]=True
    close[hanger_375,doorjamb_347]=True
    close[hanger_375,dresser_358]=True
    close[hanger_375,hanger_359]=True
    close[hanger_375,hanger_361]=True
    close[hanger_375,hanger_363]=True
    close[hanger_375,hanger_365]=True
    close[hanger_375,hanger_367]=True
    close[hanger_375,hanger_369]=True
    close[hanger_375,hanger_372]=True
    close[hanger_375,hanger_374]=True
    close[hanger_375,hanger_376]=True
    close[hanger_375,closetdrawer_377]=True
    close[hanger_375,closetdrawer_380]=True
    close[hanger_375,closetdrawer_382]=True
    close[hanger_375,closetdrawer_384]=True
    close[hanger_375,closetdrawer_388]=True
    close[hanger_376,wall_334]=True
    close[hanger_376,wall_336]=True
    close[hanger_376,ceiling_344]=True
    close[hanger_376,ceiling_345]=True
    close[hanger_376,doorjamb_347]=True
    close[hanger_376,dresser_358]=True
    close[hanger_376,hanger_359]=True
    close[hanger_376,hanger_361]=True
    close[hanger_376,hanger_363]=True
    close[hanger_376,hanger_365]=True
    close[hanger_376,hanger_367]=True
    close[hanger_376,hanger_369]=True
    close[hanger_376,hanger_372]=True
    close[hanger_376,hanger_374]=True
    close[hanger_376,hanger_375]=True
    close[hanger_376,closetdrawer_377]=True
    close[hanger_376,closetdrawer_380]=True
    close[hanger_376,closetdrawer_382]=True
    close[hanger_376,closetdrawer_384]=True
    close[hanger_376,closetdrawer_388]=True
    close[closetdrawer_377,floor_327]=True
    close[closetdrawer_377,floor_328]=True
    close[closetdrawer_377,wall_334]=True
    close[closetdrawer_377,wall_336]=True
    close[closetdrawer_377,dresser_358]=True
    close[closetdrawer_377,hanger_359]=True
    close[closetdrawer_377,hanger_361]=True
    close[closetdrawer_377,hanger_363]=True
    close[closetdrawer_377,hanger_365]=True
    close[closetdrawer_377,hanger_367]=True
    close[closetdrawer_377,hanger_369]=True
    close[closetdrawer_377,hanger_372]=True
    close[closetdrawer_377,hanger_374]=True
    close[closetdrawer_377,hanger_375]=True
    close[closetdrawer_377,hanger_376]=True
    close[closetdrawer_377,closetdrawer_380]=True
    close[closetdrawer_377,closetdrawer_382]=True
    close[closetdrawer_377,closetdrawer_384]=True
    close[closetdrawer_377,closetdrawer_388]=True
    close[closetdrawer_377,closetdrawer_392]=True
    close[closetdrawer_377,closetdrawer_394]=True
    close[closetdrawer_380,floor_327]=True
    close[closetdrawer_380,floor_328]=True
    close[closetdrawer_380,wall_334]=True
    close[closetdrawer_380,wall_336]=True
    close[closetdrawer_380,doorjamb_347]=True
    close[closetdrawer_380,dresser_358]=True
    close[closetdrawer_380,hanger_359]=True
    close[closetdrawer_380,hanger_361]=True
    close[closetdrawer_380,hanger_363]=True
    close[closetdrawer_380,hanger_365]=True
    close[closetdrawer_380,hanger_367]=True
    close[closetdrawer_380,hanger_369]=True
    close[closetdrawer_380,hanger_372]=True
    close[closetdrawer_380,hanger_374]=True
    close[closetdrawer_380,hanger_375]=True
    close[closetdrawer_380,hanger_376]=True
    close[closetdrawer_380,closetdrawer_377]=True
    close[closetdrawer_380,closetdrawer_382]=True
    close[closetdrawer_380,closetdrawer_384]=True
    close[closetdrawer_380,closetdrawer_388]=True
    close[closetdrawer_380,closetdrawer_392]=True
    close[closetdrawer_380,closetdrawer_394]=True
    close[closetdrawer_382,floor_327]=True
    close[closetdrawer_382,floor_328]=True
    close[closetdrawer_382,wall_334]=True
    close[closetdrawer_382,wall_336]=True
    close[closetdrawer_382,doorjamb_347]=True
    close[closetdrawer_382,dresser_358]=True
    close[closetdrawer_382,hanger_359]=True
    close[closetdrawer_382,hanger_363]=True
    close[closetdrawer_382,hanger_365]=True
    close[closetdrawer_382,hanger_372]=True
    close[closetdrawer_382,hanger_374]=True
    close[closetdrawer_382,hanger_375]=True
    close[closetdrawer_382,hanger_376]=True
    close[closetdrawer_382,closetdrawer_377]=True
    close[closetdrawer_382,closetdrawer_380]=True
    close[closetdrawer_382,closetdrawer_384]=True
    close[closetdrawer_382,closetdrawer_388]=True
    close[closetdrawer_382,closetdrawer_392]=True
    close[closetdrawer_382,closetdrawer_394]=True
    close[closetdrawer_384,floor_327]=True
    close[closetdrawer_384,floor_328]=True
    close[closetdrawer_384,wall_334]=True
    close[closetdrawer_384,wall_336]=True
    close[closetdrawer_384,dresser_358]=True
    close[closetdrawer_384,hanger_359]=True
    close[closetdrawer_384,hanger_361]=True
    close[closetdrawer_384,hanger_363]=True
    close[closetdrawer_384,hanger_365]=True
    close[closetdrawer_384,hanger_367]=True
    close[closetdrawer_384,hanger_369]=True
    close[closetdrawer_384,hanger_372]=True
    close[closetdrawer_384,hanger_374]=True
    close[closetdrawer_384,hanger_375]=True
    close[closetdrawer_384,hanger_376]=True
    close[closetdrawer_384,closetdrawer_377]=True
    close[closetdrawer_384,closetdrawer_380]=True
    close[closetdrawer_384,closetdrawer_382]=True
    close[closetdrawer_384,closetdrawer_388]=True
    close[closetdrawer_384,closetdrawer_392]=True
    close[closetdrawer_384,closetdrawer_394]=True
    close[closetdrawer_388,floor_327]=True
    close[closetdrawer_388,floor_328]=True
    close[closetdrawer_388,wall_334]=True
    close[closetdrawer_388,wall_336]=True
    close[closetdrawer_388,dresser_358]=True
    close[closetdrawer_388,hanger_359]=True
    close[closetdrawer_388,hanger_361]=True
    close[closetdrawer_388,hanger_363]=True
    close[closetdrawer_388,hanger_365]=True
    close[closetdrawer_388,hanger_367]=True
    close[closetdrawer_388,hanger_369]=True
    close[closetdrawer_388,hanger_372]=True
    close[closetdrawer_388,hanger_374]=True
    close[closetdrawer_388,hanger_375]=True
    close[closetdrawer_388,hanger_376]=True
    close[closetdrawer_388,closetdrawer_377]=True
    close[closetdrawer_388,closetdrawer_380]=True
    close[closetdrawer_388,closetdrawer_382]=True
    close[closetdrawer_388,closetdrawer_384]=True
    close[closetdrawer_388,closetdrawer_392]=True
    close[closetdrawer_388,closetdrawer_394]=True
    close[closetdrawer_392,floor_327]=True
    close[closetdrawer_392,floor_328]=True
    close[closetdrawer_392,wall_334]=True
    close[closetdrawer_392,wall_336]=True
    close[closetdrawer_392,doorjamb_347]=True
    close[closetdrawer_392,dresser_358]=True
    close[closetdrawer_392,closetdrawer_377]=True
    close[closetdrawer_392,closetdrawer_380]=True
    close[closetdrawer_392,closetdrawer_382]=True
    close[closetdrawer_392,closetdrawer_384]=True
    close[closetdrawer_392,closetdrawer_388]=True
    close[closetdrawer_392,closetdrawer_394]=True
    close[closetdrawer_394,floor_327]=True
    close[closetdrawer_394,floor_328]=True
    close[closetdrawer_394,wall_334]=True
    close[closetdrawer_394,wall_336]=True
    close[closetdrawer_394,dresser_358]=True
    close[closetdrawer_394,closetdrawer_377]=True
    close[closetdrawer_394,closetdrawer_380]=True
    close[closetdrawer_394,closetdrawer_382]=True
    close[closetdrawer_394,closetdrawer_384]=True
    close[closetdrawer_394,closetdrawer_388]=True
    close[closetdrawer_394,closetdrawer_392]=True
    close[filing_cabinet_399,floor_205]=True
    close[filing_cabinet_399,floor_208]=True
    close[filing_cabinet_399,wall_213]=True
    close[filing_cabinet_399,wall_214]=True
    close[filing_cabinet_399,wallshelf_235]=True
    close[filing_cabinet_399,drawing_241]=True
    close[filing_cabinet_399,drawing_242]=True
    close[filing_cabinet_399,drawing_243]=True
    close[filing_cabinet_399,floor_320]=True
    close[filing_cabinet_399,floor_325]=True
    close[filing_cabinet_399,wall_331]=True
    close[filing_cabinet_399,wall_332]=True
    close[filing_cabinet_399,doorjamb_346]=True
    close[filing_cabinet_399,bookshelf_354]=True
    close[filing_cabinet_399,drawing_402]=True
    close[filing_cabinet_399,drawing_403]=True
    close[filing_cabinet_399,drawing_404]=True
    close[filing_cabinet_399,light_411]=True
    close[filing_cabinet_399,photoframe_430]=True
    close[drawing_400,wall_333]=True
    close[drawing_400,wall_335]=True
    close[drawing_400,ceiling_338]=True
    close[drawing_400,ceiling_339]=True
    close[drawing_400,couch_352]=True
    close[drawing_400,mat_401]=True
    close[drawing_400,pillow_405]=True
    close[drawing_400,pillow_406]=True
    close[mat_401,floor_321]=True
    close[mat_401,floor_322]=True
    close[mat_401,floor_323]=True
    close[mat_401,floor_324]=True
    close[mat_401,wall_329]=True
    close[mat_401,wall_333]=True
    close[mat_401,wall_335]=True
    close[mat_401,window_348]=True
    close[mat_401,walllamp_350]=True
    close[mat_401,couch_352]=True
    close[mat_401,tvstand_353]=True
    close[mat_401,table_355]=True
    close[mat_401,drawing_400]=True
    close[mat_401,pillow_405]=True
    close[mat_401,pillow_406]=True
    close[mat_401,curtain_409]=True
    close[mat_401,television_410]=True
    close[drawing_402,wall_213]=True
    close[drawing_402,wall_214]=True
    close[drawing_402,ceiling_219]=True
    close[drawing_402,ceiling_220]=True
    close[drawing_402,table_226]=True
    close[drawing_402,wallshelf_235]=True
    close[drawing_402,drawing_241]=True
    close[drawing_402,drawing_242]=True
    close[drawing_402,drawing_243]=True
    close[drawing_402,wall_331]=True
    close[drawing_402,wall_332]=True
    close[drawing_402,ceiling_337]=True
    close[drawing_402,ceiling_342]=True
    close[drawing_402,doorjamb_346]=True
    close[drawing_402,bookshelf_354]=True
    close[drawing_402,filing_cabinet_399]=True
    close[drawing_402,drawing_403]=True
    close[drawing_402,drawing_404]=True
    close[drawing_402,light_411]=True
    close[drawing_403,wall_212]=True
    close[drawing_403,wall_213]=True
    close[drawing_403,wall_214]=True
    close[drawing_403,wall_215]=True
    close[drawing_403,ceiling_220]=True
    close[drawing_403,ceiling_221]=True
    close[drawing_403,table_226]=True
    close[drawing_403,wallshelf_234]=True
    close[drawing_403,wallshelf_235]=True
    close[drawing_403,drawing_241]=True
    close[drawing_403,drawing_242]=True
    close[drawing_403,drawing_243]=True
    close[drawing_403,wall_331]=True
    close[drawing_403,wall_332]=True
    close[drawing_403,ceiling_337]=True
    close[drawing_403,bookshelf_354]=True
    close[drawing_403,filing_cabinet_399]=True
    close[drawing_403,drawing_402]=True
    close[drawing_403,drawing_404]=True
    close[drawing_403,photoframe_430]=True
    close[drawing_404,wall_213]=True
    close[drawing_404,wall_214]=True
    close[drawing_404,ceiling_219]=True
    close[drawing_404,ceiling_220]=True
    close[drawing_404,wallshelf_235]=True
    close[drawing_404,drawing_241]=True
    close[drawing_404,drawing_242]=True
    close[drawing_404,drawing_243]=True
    close[drawing_404,wall_331]=True
    close[drawing_404,wall_332]=True
    close[drawing_404,ceiling_337]=True
    close[drawing_404,ceiling_342]=True
    close[drawing_404,doorjamb_346]=True
    close[drawing_404,filing_cabinet_399]=True
    close[drawing_404,drawing_402]=True
    close[drawing_404,drawing_403]=True
    close[drawing_404,light_411]=True
    close[pillow_405,floor_322]=True
    close[pillow_405,floor_323]=True
    close[pillow_405,wall_329]=True
    close[pillow_405,wall_333]=True
    close[pillow_405,window_348]=True
    close[pillow_405,couch_352]=True
    close[pillow_405,drawing_400]=True
    close[pillow_405,mat_401]=True
    close[pillow_405,curtain_409]=True
    close[pillow_406,floor_321]=True
    close[pillow_406,floor_322]=True
    close[pillow_406,wall_333]=True
    close[pillow_406,wall_335]=True
    close[pillow_406,walllamp_350]=True
    close[pillow_406,couch_352]=True
    close[pillow_406,table_355]=True
    close[pillow_406,drawing_400]=True
    close[pillow_406,mat_401]=True
    close[curtain_407,floor_323]=True
    close[curtain_407,wall_329]=True
    close[curtain_407,wall_334]=True
    close[curtain_407,ceiling_340]=True
    close[curtain_407,ceiling_345]=True
    close[curtain_407,window_348]=True
    close[curtain_407,couch_352]=True
    close[curtain_407,curtain_408]=True
    close[curtain_407,curtain_409]=True
    close[curtain_408,floor_323]=True
    close[curtain_408,wall_329]=True
    close[curtain_408,wall_334]=True
    close[curtain_408,ceiling_340]=True
    close[curtain_408,ceiling_345]=True
    close[curtain_408,window_348]=True
    close[curtain_408,couch_352]=True
    close[curtain_408,curtain_407]=True
    close[curtain_408,curtain_409]=True
    close[curtain_409,floor_323]=True
    close[curtain_409,wall_329]=True
    close[curtain_409,wall_333]=True
    close[curtain_409,ceiling_339]=True
    close[curtain_409,ceiling_340]=True
    close[curtain_409,window_348]=True
    close[curtain_409,couch_352]=True
    close[curtain_409,mat_401]=True
    close[curtain_409,pillow_405]=True
    close[curtain_409,curtain_407]=True
    close[curtain_409,curtain_408]=True
    close[television_410,floor_323]=True
    close[television_410,floor_324]=True
    close[television_410,floor_327]=True
    close[television_410,floor_328]=True
    close[television_410,wall_334]=True
    close[television_410,ceiling_340]=True
    close[television_410,ceiling_341]=True
    close[television_410,ceilinglamp_349]=True
    close[television_410,couch_352]=True
    close[television_410,tvstand_353]=True
    close[television_410,table_355]=True
    close[television_410,mat_401]=True
    close[light_411,floor_205]=True
    close[light_411,floor_208]=True
    close[light_411,wall_213]=True
    close[light_411,wall_214]=True
    close[light_411,ceiling_219]=True
    close[light_411,ceiling_220]=True
    close[light_411,wallshelf_235]=True
    close[light_411,floor_320]=True
    close[light_411,floor_325]=True
    close[light_411,wall_331]=True
    close[light_411,wall_332]=True
    close[light_411,ceiling_337]=True
    close[light_411,ceiling_342]=True
    close[light_411,doorjamb_346]=True
    close[light_411,filing_cabinet_399]=True
    close[light_411,drawing_402]=True
    close[light_411,drawing_404]=True
    close[powersocket_412,floor_208]=True
    close[powersocket_412,wall_213]=True
    close[powersocket_412,tvstand_225]=True
    close[powersocket_412,floor_325]=True
    close[powersocket_412,floor_326]=True
    close[powersocket_412,wall_330]=True
    close[powersocket_412,wall_331]=True
    close[powersocket_412,doorjamb_346]=True
    close[powersocket_412,desk_357]=True
    close[powersocket_412,mouse_413]=True
    close[powersocket_412,mousepad_414]=True
    close[powersocket_412,computer_417]=True
    close[mouse_413,floor_208]=True
    close[mouse_413,wall_213]=True
    close[mouse_413,floor_325]=True
    close[mouse_413,floor_326]=True
    close[mouse_413,wall_330]=True
    close[mouse_413,wall_331]=True
    close[mouse_413,doorjamb_346]=True
    close[mouse_413,chair_356]=True
    close[mouse_413,desk_357]=True
    close[mouse_413,powersocket_412]=True
    close[mouse_413,mousepad_414]=True
    close[mouse_413,keyboard_415]=True
    close[mouse_413,cpuscreen_416]=True
    close[mouse_413,computer_417]=True
    close[mousepad_414,floor_208]=True
    close[mousepad_414,wall_213]=True
    close[mousepad_414,floor_325]=True
    close[mousepad_414,floor_326]=True
    close[mousepad_414,wall_330]=True
    close[mousepad_414,wall_331]=True
    close[mousepad_414,doorjamb_346]=True
    close[mousepad_414,chair_356]=True
    close[mousepad_414,desk_357]=True
    close[mousepad_414,powersocket_412]=True
    close[mousepad_414,mouse_413]=True
    close[mousepad_414,keyboard_415]=True
    close[mousepad_414,cpuscreen_416]=True
    close[mousepad_414,computer_417]=True
    close[keyboard_415,wall_213]=True
    close[keyboard_415,floor_325]=True
    close[keyboard_415,floor_326]=True
    close[keyboard_415,wall_330]=True
    close[keyboard_415,wall_331]=True
    close[keyboard_415,walllamp_351]=True
    close[keyboard_415,chair_356]=True
    close[keyboard_415,desk_357]=True
    close[keyboard_415,mouse_413]=True
    close[keyboard_415,mousepad_414]=True
    close[keyboard_415,cpuscreen_416]=True
    close[keyboard_415,computer_417]=True
    close[cpuscreen_416,wall_213]=True
    close[cpuscreen_416,floor_326]=True
    close[cpuscreen_416,wall_330]=True
    close[cpuscreen_416,wall_331]=True
    close[cpuscreen_416,ceiling_343]=True
    close[cpuscreen_416,chair_356]=True
    close[cpuscreen_416,desk_357]=True
    close[cpuscreen_416,mouse_413]=True
    close[cpuscreen_416,mousepad_414]=True
    close[cpuscreen_416,keyboard_415]=True
    close[cpuscreen_416,computer_417]=True
    close[computer_417,floor_208]=True
    close[computer_417,wall_213]=True
    close[computer_417,floor_325]=True
    close[computer_417,floor_326]=True
    close[computer_417,wall_330]=True
    close[computer_417,wall_331]=True
    close[computer_417,doorjamb_346]=True
    close[computer_417,chair_356]=True
    close[computer_417,desk_357]=True
    close[computer_417,powersocket_412]=True
    close[computer_417,mouse_413]=True
    close[computer_417,mousepad_414]=True
    close[computer_417,keyboard_415]=True
    close[computer_417,cpuscreen_416]=True
    close[photoframe_430,wall_212]=True
    close[photoframe_430,wall_214]=True
    close[photoframe_430,wall_215]=True
    close[photoframe_430,wallshelf_234]=True
    close[photoframe_430,drawing_241]=True
    close[photoframe_430,drawing_243]=True
    close[photoframe_430,floor_320]=True
    close[photoframe_430,wall_332]=True
    close[photoframe_430,wall_335]=True
    close[photoframe_430,ceiling_337]=True
    close[photoframe_430,bookshelf_354]=True
    close[photoframe_430,filing_cabinet_399]=True
    close[photoframe_430,drawing_403]=True
    close[plate_1000,sink_231]=True
    close[dishwasher_1001,sink_231]=True
    close[coffee_filter_2000,table_226]=True
    close[pencil_2001,desk_357]=True
    close[hairbrush_2002,couch_352]=True
    close[drawing_2003,table_226]=True
    close[chair_2004,floor_69]=True
    close[napkin_2005,kitchen_counter_230]=True
    facing[floor_2,drawing_174]=True
    facing[floor_3,drawing_174]=True
    facing[floor_6,drawing_174]=True
    facing[wall_12,drawing_174]=True
    facing[wall_14,drawing_174]=True
    facing[ceiling_16,drawing_174]=True
    facing[ceiling_17,drawing_174]=True
    facing[mat_22,drawing_174]=True
    facing[door_44,drawing_174]=True
    facing[doorjamb_45,drawing_174]=True
    facing[floor_68,drawing_175]=True
    facing[floor_69,drawing_175]=True
    facing[floor_70,drawing_176]=True
    facing[floor_71,drawing_176]=True
    facing[floor_72,computer_170]=True
    facing[floor_72,drawing_174]=True
    facing[floor_72,drawing_176]=True
    facing[floor_73,computer_170]=True
    facing[floor_73,drawing_174]=True
    facing[floor_73,drawing_175]=True
    facing[floor_73,drawing_176]=True
    facing[floor_74,computer_170]=True
    facing[floor_74,drawing_175]=True
    facing[floor_75,computer_170]=True
    facing[floor_75,drawing_175]=True
    facing[floor_76,computer_170]=True
    facing[floor_76,drawing_174]=True
    facing[floor_76,drawing_175]=True
    facing[floor_77,drawing_174]=True
    facing[wall_78,computer_170]=True
    facing[wall_79,drawing_174]=True
    facing[wall_80,drawing_176]=True
    facing[wall_81,drawing_175]=True
    facing[wall_82,drawing_176]=True
    facing[wall_83,computer_170]=True
    facing[wall_83,drawing_175]=True
    facing[wall_84,drawing_175]=True
    facing[wall_84,drawing_242]=True
    facing[wall_85,drawing_174]=True
    facing[window_86,drawing_176]=True
    facing[ceiling_87,drawing_175]=True
    facing[ceiling_88,drawing_176]=True
    facing[ceiling_89,drawing_176]=True
    facing[ceiling_90,drawing_174]=True
    facing[ceiling_90,drawing_176]=True
    facing[ceiling_91,computer_170]=True
    facing[ceiling_91,drawing_174]=True
    facing[ceiling_91,drawing_175]=True
    facing[ceiling_91,drawing_176]=True
    facing[ceiling_92,computer_170]=True
    facing[ceiling_92,drawing_175]=True
    facing[ceiling_93,computer_170]=True
    facing[ceiling_93,drawing_175]=True
    facing[ceiling_94,computer_170]=True
    facing[ceiling_94,drawing_174]=True
    facing[ceiling_94,drawing_175]=True
    facing[ceiling_95,drawing_174]=True
    facing[ceilinglamp_96,computer_170]=True
    facing[ceilinglamp_96,drawing_174]=True
    facing[ceilinglamp_96,drawing_175]=True
    facing[ceilinglamp_96,drawing_176]=True
    facing[tablelamp_98,drawing_176]=True
    facing[trashcan_99,drawing_238]=True
    facing[trashcan_99,drawing_239]=True
    facing[trashcan_99,drawing_240]=True
    facing[trashcan_99,drawing_243]=True
    facing[bookshelf_101,drawing_174]=True
    facing[nightstand_102,drawing_176]=True
    facing[desk_104,drawing_175]=True
    facing[bed_105,drawing_176]=True
    facing[chair_106,drawing_176]=True
    facing[table_107,computer_170]=True
    facing[table_107,drawing_174]=True
    facing[table_107,drawing_175]=True
    facing[table_107,drawing_176]=True
    facing[dresser_108,computer_170]=True
    facing[hanger_112,computer_170]=True
    facing[hanger_113,computer_170]=True
    facing[hanger_115,computer_170]=True
    facing[doorjamb_165,drawing_242]=True
    facing[doorjamb_165,drawing_243]=True
    facing[doorjamb_165,wall_clock_249]=True
    facing[mouse_166,drawing_175]=True
    facing[mousepad_167,drawing_175]=True
    facing[keyboard_168,drawing_175]=True
    facing[light_169,drawing_175]=True
    facing[cpuscreen_171,drawing_175]=True
    facing[mat_173,drawing_176]=True
    facing[orchid_178,computer_170]=True
    facing[orchid_178,drawing_174]=True
    facing[orchid_178,drawing_175]=True
    facing[orchid_178,drawing_176]=True
    facing[curtain_179,drawing_176]=True
    facing[curtain_180,drawing_176]=True
    facing[curtain_181,drawing_176]=True
    facing[pillow_182,drawing_176]=True
    facing[pillow_183,drawing_176]=True
    facing[photoframe_185,drawing_174]=True
    facing[floor_202,drawing_238]=True
    facing[floor_202,drawing_239]=True
    facing[floor_202,drawing_240]=True
    facing[floor_202,drawing_241]=True
    facing[floor_202,drawing_242]=True
    facing[floor_202,drawing_243]=True
    facing[floor_203,drawing_238]=True
    facing[floor_203,drawing_239]=True
    facing[floor_203,drawing_240]=True
    facing[floor_203,drawing_241]=True
    facing[floor_203,drawing_242]=True
    facing[floor_203,drawing_243]=True
    facing[floor_204,drawing_238]=True
    facing[floor_204,drawing_239]=True
    facing[floor_204,drawing_240]=True
    facing[floor_204,drawing_241]=True
    facing[floor_204,drawing_242]=True
    facing[floor_204,drawing_243]=True
    facing[floor_205,drawing_238]=True
    facing[floor_205,drawing_239]=True
    facing[floor_205,drawing_240]=True
    facing[floor_205,drawing_241]=True
    facing[floor_205,drawing_242]=True
    facing[floor_205,drawing_243]=True
    facing[floor_206,drawing_238]=True
    facing[floor_206,drawing_239]=True
    facing[floor_206,drawing_240]=True
    facing[floor_206,drawing_241]=True
    facing[floor_206,drawing_242]=True
    facing[floor_206,drawing_243]=True
    facing[floor_206,television_248]=True
    facing[floor_206,wall_clock_249]=True
    facing[floor_207,drawing_238]=True
    facing[floor_207,drawing_240]=True
    facing[floor_207,drawing_242]=True
    facing[floor_207,drawing_243]=True
    facing[floor_207,television_248]=True
    facing[floor_208,drawing_241]=True
    facing[floor_208,drawing_242]=True
    facing[floor_208,drawing_243]=True
    facing[wall_209,drawing_241]=True
    facing[wall_209,drawing_242]=True
    facing[wall_209,drawing_243]=True
    facing[wall_209,television_248]=True
    facing[wall_209,wall_clock_249]=True
    facing[wall_210,drawing_238]=True
    facing[wall_210,drawing_240]=True
    facing[wall_210,drawing_241]=True
    facing[wall_210,drawing_242]=True
    facing[wall_210,drawing_243]=True
    facing[wall_210,television_248]=True
    facing[wall_210,wall_clock_249]=True
    facing[wall_211,drawing_238]=True
    facing[wall_211,drawing_239]=True
    facing[wall_211,drawing_240]=True
    facing[wall_211,drawing_241]=True
    facing[wall_211,drawing_242]=True
    facing[wall_211,drawing_243]=True
    facing[wall_212,drawing_238]=True
    facing[wall_212,drawing_239]=True
    facing[wall_212,drawing_240]=True
    facing[wall_212,drawing_241]=True
    facing[wall_212,drawing_242]=True
    facing[wall_212,drawing_243]=True
    facing[wall_213,drawing_241]=True
    facing[wall_213,drawing_242]=True
    facing[wall_213,drawing_243]=True
    facing[wall_213,television_248]=True
    facing[wall_214,television_248]=True
    facing[wall_215,drawing_404]=True
    facing[ceiling_216,drawing_238]=True
    facing[ceiling_216,drawing_239]=True
    facing[ceiling_216,drawing_240]=True
    facing[ceiling_216,drawing_241]=True
    facing[ceiling_216,drawing_242]=True
    facing[ceiling_216,drawing_243]=True
    facing[ceiling_217,drawing_238]=True
    facing[ceiling_217,drawing_239]=True
    facing[ceiling_217,drawing_240]=True
    facing[ceiling_217,drawing_241]=True
    facing[ceiling_217,drawing_242]=True
    facing[ceiling_217,drawing_243]=True
    facing[ceiling_217,television_248]=True
    facing[ceiling_217,wall_clock_249]=True
    facing[ceiling_218,drawing_238]=True
    facing[ceiling_218,drawing_240]=True
    facing[ceiling_218,drawing_241]=True
    facing[ceiling_218,drawing_242]=True
    facing[ceiling_218,television_248]=True
    facing[ceiling_218,wall_clock_249]=True
    facing[ceiling_219,drawing_241]=True
    facing[ceiling_219,drawing_242]=True
    facing[ceiling_219,drawing_243]=True
    facing[ceiling_219,television_248]=True
    facing[ceiling_220,drawing_238]=True
    facing[ceiling_220,drawing_239]=True
    facing[ceiling_220,drawing_240]=True
    facing[ceiling_220,drawing_241]=True
    facing[ceiling_220,drawing_242]=True
    facing[ceiling_220,drawing_243]=True
    facing[ceiling_220,television_248]=True
    facing[ceiling_221,drawing_238]=True
    facing[ceiling_221,drawing_239]=True
    facing[ceiling_221,drawing_240]=True
    facing[ceiling_221,drawing_241]=True
    facing[ceiling_221,drawing_242]=True
    facing[ceiling_221,drawing_243]=True
    facing[door_222,television_248]=True
    facing[door_222,wall_clock_249]=True
    facing[ceilinglamp_223,drawing_238]=True
    facing[ceilinglamp_223,drawing_239]=True
    facing[ceilinglamp_223,drawing_240]=True
    facing[ceilinglamp_223,drawing_241]=True
    facing[ceilinglamp_223,drawing_242]=True
    facing[ceilinglamp_223,drawing_243]=True
    facing[ceilinglamp_223,television_248]=True
    facing[ceilinglamp_223,wall_clock_249]=True
    facing[ceilinglamp_224,drawing_238]=True
    facing[ceilinglamp_224,drawing_239]=True
    facing[ceilinglamp_224,drawing_240]=True
    facing[ceilinglamp_224,drawing_241]=True
    facing[ceilinglamp_224,drawing_242]=True
    facing[ceilinglamp_224,drawing_243]=True
    facing[ceilinglamp_224,television_248]=True
    facing[tvstand_225,drawing_241]=True
    facing[tvstand_225,drawing_242]=True
    facing[tvstand_225,drawing_243]=True
    facing[table_226,drawing_238]=True
    facing[table_226,drawing_239]=True
    facing[table_226,drawing_240]=True
    facing[table_226,drawing_241]=True
    facing[table_226,drawing_242]=True
    facing[table_226,drawing_243]=True
    facing[table_226,television_248]=True
    facing[bench_227,drawing_238]=True
    facing[bench_227,drawing_239]=True
    facing[bench_227,drawing_240]=True
    facing[bench_227,drawing_241]=True
    facing[bench_227,drawing_242]=True
    facing[bench_227,drawing_243]=True
    facing[bench_227,television_248]=True
    facing[bench_227,wall_clock_249]=True
    facing[bench_228,drawing_238]=True
    facing[bench_228,drawing_239]=True
    facing[bench_228,drawing_240]=True
    facing[bench_228,drawing_241]=True
    facing[bench_228,drawing_242]=True
    facing[bench_228,drawing_243]=True
    facing[kitchen_counter_230,drawing_238]=True
    facing[kitchen_counter_230,drawing_239]=True
    facing[kitchen_counter_230,drawing_240]=True
    facing[kitchen_counter_230,drawing_241]=True
    facing[kitchen_counter_230,drawing_242]=True
    facing[kitchen_counter_230,drawing_243]=True
    facing[faucet_232,drawing_238]=True
    facing[faucet_232,drawing_239]=True
    facing[faucet_232,drawing_240]=True
    facing[faucet_232,drawing_241]=True
    facing[faucet_232,drawing_242]=True
    facing[faucet_232,drawing_243]=True
    facing[bookshelf_233,television_248]=True
    facing[wallshelf_234,drawing_238]=True
    facing[wallshelf_234,drawing_239]=True
    facing[wallshelf_234,drawing_240]=True
    facing[wallshelf_235,television_248]=True
    facing[mat_236,drawing_238]=True
    facing[mat_236,drawing_239]=True
    facing[mat_236,drawing_240]=True
    facing[mat_236,drawing_241]=True
    facing[mat_236,drawing_242]=True
    facing[mat_236,drawing_243]=True
    facing[mat_236,television_248]=True
    facing[mat_236,wall_clock_249]=True
    facing[mat_237,drawing_238]=True
    facing[mat_237,drawing_239]=True
    facing[mat_237,drawing_240]=True
    facing[mat_237,drawing_241]=True
    facing[mat_237,drawing_242]=True
    facing[mat_237,drawing_243]=True
    facing[mat_237,wall_clock_249]=True
    facing[drawing_238,drawing_241]=True
    facing[drawing_238,drawing_243]=True
    facing[drawing_241,drawing_238]=True
    facing[drawing_241,television_248]=True
    facing[drawing_242,television_248]=True
    facing[drawing_243,drawing_238]=True
    facing[drawing_243,television_248]=True
    facing[orchid_244,drawing_241]=True
    facing[orchid_244,drawing_242]=True
    facing[orchid_244,drawing_243]=True
    facing[orchid_244,television_248]=True
    facing[light_245,drawing_241]=True
    facing[light_245,drawing_242]=True
    facing[light_245,drawing_243]=True
    facing[light_245,television_248]=True
    facing[light_245,wall_clock_249]=True
    facing[powersocket_246,drawing_243]=True
    facing[powersocket_246,wall_clock_249]=True
    facing[phone_247,drawing_241]=True
    facing[phone_247,drawing_242]=True
    facing[phone_247,drawing_243]=True
    facing[phone_247,television_248]=True
    facing[phone_247,wall_clock_249]=True
    facing[television_248,drawing_241]=True
    facing[television_248,drawing_242]=True
    facing[television_248,drawing_243]=True
    facing[television_248,wall_clock_249]=True
    facing[wall_clock_249,drawing_241]=True
    facing[wall_clock_249,drawing_242]=True
    facing[wall_clock_249,drawing_243]=True
    facing[wall_clock_249,television_248]=True
    facing[photoframe_285,drawing_241]=True
    facing[photoframe_285,drawing_242]=True
    facing[photoframe_285,drawing_243]=True
    facing[stovefan_288,drawing_238]=True
    facing[stovefan_288,drawing_239]=True
    facing[stovefan_288,drawing_240]=True
    facing[fridge_289,drawing_239]=True
    facing[coffe_maker_290,drawing_238]=True
    facing[coffe_maker_290,drawing_239]=True
    facing[coffe_maker_290,drawing_240]=True
    facing[coffe_maker_290,drawing_241]=True
    facing[coffe_maker_290,drawing_242]=True
    facing[coffe_maker_290,drawing_243]=True
    facing[toaster_292,drawing_238]=True
    facing[toaster_292,drawing_239]=True
    facing[toaster_292,drawing_240]=True
    facing[toaster_292,drawing_241]=True
    facing[toaster_292,drawing_242]=True
    facing[toaster_292,drawing_243]=True
    facing[oven_295,drawing_238]=True
    facing[oven_295,drawing_239]=True
    facing[oven_295,drawing_240]=True
    facing[microwave_297,drawing_238]=True
    facing[microwave_297,drawing_239]=True
    facing[microwave_297,drawing_240]=True
    facing[microwave_297,drawing_241]=True
    facing[microwave_297,drawing_242]=True
    facing[microwave_297,drawing_243]=True
    facing[floor_320,drawing_400]=True
    facing[floor_320,drawing_402]=True
    facing[floor_320,drawing_403]=True
    facing[floor_320,drawing_404]=True
    facing[floor_320,television_410]=True
    facing[floor_321,drawing_400]=True
    facing[floor_321,drawing_402]=True
    facing[floor_321,drawing_403]=True
    facing[floor_321,drawing_404]=True
    facing[floor_323,drawing_400]=True
    facing[floor_324,drawing_400]=True
    facing[floor_324,drawing_402]=True
    facing[floor_324,drawing_403]=True
    facing[floor_324,drawing_404]=True
    facing[floor_324,television_410]=True
    facing[floor_324,computer_417]=True
    facing[floor_325,drawing_402]=True
    facing[floor_325,drawing_403]=True
    facing[floor_325,drawing_404]=True
    facing[floor_326,drawing_402]=True
    facing[floor_326,drawing_404]=True
    facing[floor_326,computer_417]=True
    facing[floor_327,computer_417]=True
    facing[wall_329,drawing_400]=True
    facing[wall_330,drawing_402]=True
    facing[wall_330,drawing_404]=True
    facing[wall_330,computer_417]=True
    facing[wall_332,drawing_400]=True
    facing[wall_332,drawing_402]=True
    facing[wall_332,drawing_403]=True
    facing[wall_332,drawing_404]=True
    facing[wall_332,television_410]=True
    facing[wall_333,drawing_400]=True
    facing[wall_333,television_410]=True
    facing[wall_335,drawing_402]=True
    facing[wall_335,drawing_403]=True
    facing[wall_335,drawing_404]=True
    facing[wall_335,television_410]=True
    facing[wall_336,computer_417]=True
    facing[ceiling_337,drawing_400]=True
    facing[ceiling_337,drawing_402]=True
    facing[ceiling_337,drawing_403]=True
    facing[ceiling_337,drawing_404]=True
    facing[ceiling_338,drawing_400]=True
    facing[ceiling_338,drawing_402]=True
    facing[ceiling_338,drawing_403]=True
    facing[ceiling_338,drawing_404]=True
    facing[ceiling_338,television_410]=True
    facing[ceiling_339,drawing_400]=True
    facing[ceiling_339,television_410]=True
    facing[ceiling_340,drawing_400]=True
    facing[ceiling_340,television_410]=True
    facing[ceiling_341,drawing_400]=True
    facing[ceiling_341,drawing_402]=True
    facing[ceiling_341,drawing_403]=True
    facing[ceiling_341,drawing_404]=True
    facing[ceiling_341,television_410]=True
    facing[ceiling_341,computer_417]=True
    facing[ceiling_342,drawing_402]=True
    facing[ceiling_342,drawing_403]=True
    facing[ceiling_342,drawing_404]=True
    facing[ceiling_343,drawing_402]=True
    facing[ceiling_343,drawing_404]=True
    facing[ceiling_343,computer_417]=True
    facing[ceiling_344,computer_417]=True
    facing[doorjamb_346,television_248]=True
    facing[doorjamb_347,computer_417]=True
    facing[window_348,drawing_400]=True
    facing[ceilinglamp_349,drawing_400]=True
    facing[ceilinglamp_349,drawing_402]=True
    facing[ceilinglamp_349,drawing_403]=True
    facing[ceilinglamp_349,drawing_404]=True
    facing[ceilinglamp_349,television_410]=True
    facing[ceilinglamp_349,computer_417]=True
    facing[walllamp_350,drawing_402]=True
    facing[walllamp_350,drawing_404]=True
    facing[walllamp_350,television_410]=True
    facing[walllamp_351,computer_417]=True
    facing[couch_352,television_410]=True
    facing[tvstand_353,drawing_400]=True
    facing[tvstand_353,television_410]=True
    facing[tvstand_353,computer_417]=True
    facing[bookshelf_354,drawing_402]=True
    facing[bookshelf_354,drawing_403]=True
    facing[bookshelf_354,drawing_404]=True
    facing[table_355,drawing_400]=True
    facing[table_355,drawing_404]=True
    facing[table_355,television_410]=True
    facing[table_355,computer_417]=True
    facing[chair_356,computer_417]=True
    facing[filing_cabinet_399,drawing_402]=True
    facing[filing_cabinet_399,drawing_403]=True
    facing[filing_cabinet_399,drawing_404]=True
    facing[drawing_400,television_410]=True
    facing[mat_401,drawing_400]=True
    facing[pillow_405,drawing_400]=True
    facing[pillow_405,television_410]=True
    facing[pillow_406,drawing_400]=True
    facing[pillow_406,drawing_402]=True
    facing[pillow_406,drawing_403]=True
    facing[pillow_406,drawing_404]=True
    facing[pillow_406,television_410]=True
    facing[curtain_407,drawing_400]=True
    facing[curtain_408,drawing_400]=True
    facing[curtain_409,drawing_400]=True
    facing[curtain_409,television_410]=True
    facing[television_410,drawing_400]=True
    facing[television_410,computer_417]=True
    facing[photoframe_430,drawing_402]=True
    facing[photoframe_430,drawing_403]=True
    facing[photoframe_430,drawing_404]=True
    #relations_end

    #exploration
    #exploration_end

    #id
    id[clothes_pants_2085]=2085
    id[clothes_shirt_2086]=2086
    id[clothes_socks_2087]=2087
    id[clothes_skirt_2088]=2088
    id[iron_2089]=2089
    id[basket_for_clothes_2006]=2006
    id[washing_machine_2007]=2007
    id[food_steak_2008]=2008
    id[food_apple_2009]=2009
    id[food_bacon_2010]=2010
    id[food_banana_2011]=2011
    id[food_bread_2012]=2012
    id[food_cake_2013]=2013
    id[food_carrot_2014]=2014
    id[food_cereal_2015]=2015
    id[food_cheese_2016]=2016
    id[food_chicken_2017]=2017
    id[food_dessert_2018]=2018
    id[food_donut_2019]=2019
    id[food_egg_2020]=2020
    id[food_fish_2021]=2021
    id[food_food_2022]=2022
    id[food_fruit_2023]=2023
    id[food_hamburger_2024]=2024
    id[food_ice_cream_2025]=2025
    id[food_jam_2026]=2026
    id[food_kiwi_2027]=2027
    id[food_lemon_2028]=2028
    id[food_noodles_2029]=2029
    id[food_oatmeal_2030]=2030
    id[food_orange_2031]=2031
    id[food_onion_2032]=2032
    id[food_peanut_butter_2033]=2033
    id[food_pizza_2034]=2034
    id[food_potato_2035]=2035
    id[food_rice_2036]=2036
    id[food_salt_2037]=2037
    id[food_snack_2038]=2038
    id[food_sugar_2039]=2039
    id[food_turkey_2040]=2040
    id[food_vegetable_2041]=2041
    id[dry_pasta_2042]=2042
    id[milk_2043]=2043
    id[clothes_dress_2044]=2044
    id[clothes_hat_2045]=2045
    id[clothes_gloves_2046]=2046
    id[clothes_jacket_2047]=2047
    id[clothes_scarf_2048]=2048
    id[clothes_underwear_2049]=2049
    id[knife_2050]=2050
    id[cutting_board_2051]=2051
    id[remote_control_2052]=2052
    id[soap_2053]=2053
    id[soap_2054]=2054
    id[cat_2055]=2055
    id[towel_2056]=2056
    id[towel_2057]=2057
    id[towel_2058]=2058
    id[towel_2059]=2059
    id[cd_player_2060]=2060
    id[dvd_player_2061]=2061
    id[headset_2062]=2062
    id[cup_2063]=2063
    id[cup_2064]=2064
    id[stove_2065]=2065
    id[book_2066]=2066
    id[book_2067]=2067
    id[coffee_table_2068]=2068
    id[pot_2069]=2069
    id[vacuum_cleaner_2070]=2070
    id[bowl_2071]=2071
    id[bowl_2072]=2072
    id[cleaning_solution_2073]=2073
    id[ironing_board_2074]=2074
    id[cd_2075]=2075
    id[headset_2076]=2076
    id[phone_2077]=2077
    id[sauce_2078]=2078
    id[oil_2079]=2079
    id[fork_2080]=2080
    id[fork_2081]=2081
    id[spectacles_2082]=2082
    id[fryingpan_2083]=2083
    id[detergent_2084]=2084
    id[bathroom_1]=1
    id[floor_2]=2
    id[floor_3]=3
    id[floor_4]=4
    id[floor_5]=5
    id[floor_6]=6
    id[floor_7]=7
    id[floor_8]=8
    id[wall_9]=9
    id[wall_10]=10
    id[wall_11]=11
    id[wall_12]=12
    id[wall_13]=13
    id[wall_14]=14
    id[wall_15]=15
    id[ceiling_16]=16
    id[ceiling_17]=17
    id[ceiling_18]=18
    id[ceiling_19]=19
    id[ceiling_20]=20
    id[ceiling_21]=21
    id[mat_22]=22
    id[curtain_23]=23
    id[curtain_24]=24
    id[curtain_25]=25
    id[ceilinglamp_26]=26
    id[walllamp_27]=27
    id[walllamp_28]=28
    id[walllamp_29]=29
    id[bathtub_30]=30
    id[towel_rack_31]=31
    id[towel_rack_32]=32
    id[towel_rack_33]=33
    id[towel_rack_34]=34
    id[wallshelf_35]=35
    id[shower_36]=36
    id[toilet_37]=37
    id[shower_38]=38
    id[curtain_39]=39
    id[bathroom_cabinet_40]=40
    id[bathroom_counter_41]=41
    id[sink_42]=42
    id[faucet_43]=43
    id[door_44]=44
    id[doorjamb_45]=45
    id[window_63]=63
    id[light_64]=64
    id[bedroom_67]=67
    id[floor_68]=68
    id[floor_69]=69
    id[floor_70]=70
    id[floor_71]=71
    id[floor_72]=72
    id[floor_73]=73
    id[floor_74]=74
    id[floor_75]=75
    id[floor_76]=76
    id[floor_77]=77
    id[wall_78]=78
    id[wall_79]=79
    id[wall_80]=80
    id[wall_81]=81
    id[wall_82]=82
    id[wall_83]=83
    id[wall_84]=84
    id[wall_85]=85
    id[window_86]=86
    id[ceiling_87]=87
    id[ceiling_88]=88
    id[ceiling_89]=89
    id[ceiling_90]=90
    id[ceiling_91]=91
    id[ceiling_92]=92
    id[ceiling_93]=93
    id[ceiling_94]=94
    id[ceiling_95]=95
    id[ceilinglamp_96]=96
    id[tablelamp_97]=97
    id[tablelamp_98]=98
    id[trashcan_99]=99
    id[nightstand_100]=100
    id[bookshelf_101]=101
    id[nightstand_102]=102
    id[chair_103]=103
    id[desk_104]=104
    id[bed_105]=105
    id[chair_106]=106
    id[table_107]=107
    id[dresser_108]=108
    id[hanger_109]=109
    id[hanger_110]=110
    id[hanger_111]=111
    id[hanger_112]=112
    id[hanger_113]=113
    id[hanger_114]=114
    id[hanger_115]=115
    id[closetdrawer_116]=116
    id[closetdrawer_117]=117
    id[closetdrawer_118]=118
    id[closetdrawer_119]=119
    id[closetdrawer_120]=120
    id[closetdrawer_121]=121
    id[closetdrawer_122]=122
    id[dresser_123]=123
    id[hanger_124]=124
    id[hanger_126]=126
    id[hanger_128]=128
    id[hanger_130]=130
    id[hanger_132]=132
    id[hanger_134]=134
    id[hanger_136]=136
    id[hanger_138]=138
    id[hanger_140]=140
    id[hanger_141]=141
    id[hanger_142]=142
    id[closetdrawer_143]=143
    id[closetdrawer_146]=146
    id[closetdrawer_148]=148
    id[closetdrawer_150]=150
    id[closetdrawer_154]=154
    id[closetdrawer_158]=158
    id[closetdrawer_160]=160
    id[doorjamb_165]=165
    id[mouse_166]=166
    id[mousepad_167]=167
    id[keyboard_168]=168
    id[light_169]=169
    id[computer_170]=170
    id[cpuscreen_171]=171
    id[mat_173]=173
    id[drawing_174]=174
    id[drawing_175]=175
    id[drawing_176]=176
    id[orchid_178]=178
    id[curtain_179]=179
    id[curtain_180]=180
    id[curtain_181]=181
    id[pillow_182]=182
    id[pillow_183]=183
    id[photoframe_185]=185
    id[dining_room_201]=201
    id[floor_202]=202
    id[floor_203]=203
    id[floor_204]=204
    id[floor_205]=205
    id[floor_206]=206
    id[floor_207]=207
    id[floor_208]=208
    id[wall_209]=209
    id[wall_210]=210
    id[wall_211]=211
    id[wall_212]=212
    id[wall_213]=213
    id[wall_214]=214
    id[wall_215]=215
    id[ceiling_216]=216
    id[ceiling_217]=217
    id[ceiling_218]=218
    id[ceiling_219]=219
    id[ceiling_220]=220
    id[ceiling_221]=221
    id[door_222]=222
    id[ceilinglamp_223]=223
    id[ceilinglamp_224]=224
    id[tvstand_225]=225
    id[table_226]=226
    id[bench_227]=227
    id[bench_228]=228
    id[cupboard_229]=229
    id[kitchen_counter_230]=230
    id[sink_231]=231
    id[faucet_232]=232
    id[bookshelf_233]=233
    id[wallshelf_234]=234
    id[wallshelf_235]=235
    id[mat_236]=236
    id[mat_237]=237
    id[drawing_238]=238
    id[drawing_239]=239
    id[drawing_240]=240
    id[drawing_241]=241
    id[drawing_242]=242
    id[drawing_243]=243
    id[orchid_244]=244
    id[light_245]=245
    id[powersocket_246]=246
    id[phone_247]=247
    id[television_248]=248
    id[wall_clock_249]=249
    id[photoframe_285]=285
    id[stovefan_288]=288
    id[fridge_289]=289
    id[coffe_maker_290]=290
    id[toaster_292]=292
    id[oven_295]=295
    id[tray_296]=296
    id[microwave_297]=297
    id[home_office_319]=319
    id[floor_320]=320
    id[floor_321]=321
    id[floor_322]=322
    id[floor_323]=323
    id[floor_324]=324
    id[floor_325]=325
    id[floor_326]=326
    id[floor_327]=327
    id[floor_328]=328
    id[wall_329]=329
    id[wall_330]=330
    id[wall_331]=331
    id[wall_332]=332
    id[wall_333]=333
    id[wall_334]=334
    id[wall_335]=335
    id[wall_336]=336
    id[ceiling_337]=337
    id[ceiling_338]=338
    id[ceiling_339]=339
    id[ceiling_340]=340
    id[ceiling_341]=341
    id[ceiling_342]=342
    id[ceiling_343]=343
    id[ceiling_344]=344
    id[ceiling_345]=345
    id[doorjamb_346]=346
    id[doorjamb_347]=347
    id[window_348]=348
    id[ceilinglamp_349]=349
    id[walllamp_350]=350
    id[walllamp_351]=351
    id[couch_352]=352
    id[tvstand_353]=353
    id[bookshelf_354]=354
    id[table_355]=355
    id[chair_356]=356
    id[desk_357]=357
    id[dresser_358]=358
    id[hanger_359]=359
    id[hanger_361]=361
    id[hanger_363]=363
    id[hanger_365]=365
    id[hanger_367]=367
    id[hanger_369]=369
    id[hanger_372]=372
    id[hanger_374]=374
    id[hanger_375]=375
    id[hanger_376]=376
    id[closetdrawer_377]=377
    id[closetdrawer_380]=380
    id[closetdrawer_382]=382
    id[closetdrawer_384]=384
    id[closetdrawer_388]=388
    id[closetdrawer_392]=392
    id[closetdrawer_394]=394
    id[filing_cabinet_399]=399
    id[drawing_400]=400
    id[mat_401]=401
    id[drawing_402]=402
    id[drawing_403]=403
    id[drawing_404]=404
    id[pillow_405]=405
    id[pillow_406]=406
    id[curtain_407]=407
    id[curtain_408]=408
    id[curtain_409]=409
    id[television_410]=410
    id[light_411]=411
    id[powersocket_412]=412
    id[mouse_413]=413
    id[mousepad_414]=414
    id[keyboard_415]=415
    id[cpuscreen_416]=416
    id[computer_417]=417
    id[photoframe_430]=430
    id[plate_1000]=1000
    id[dishwasher_1001]=1001
    id[coffee_filter_2000]=2000
    id[pencil_2001]=2001
    id[hairbrush_2002]=2002
    id[drawing_2003]=2003
    id[chair_2004]=2004
    id[napkin_2005]=2005
    #id_end

    #size
    size[cup_2063]=10
    size[cup_2064]=6
    size[coffe_maker_290]=8
    #size_end
