problem "agent-problem"
domain "virtualhome_partial.cdl"

#!pragma planner_is_goal_serializable=False
#!pragma planner_is_goal_ordered=True
#!pragma planner_always_commit_skeleton=True

objects:
#objects
  keyboard_2111:item
  mouse_2112:item
  clothes_pants_2113:item
  clothes_shirt_2114:item
  clothes_socks_2115:item
  clothes_skirt_2116:item
  iron_2117:item
  chair_2118:item
  basket_for_clothes_2040:item
  washing_machine_2041:item
  food_steak_2042:item
  food_apple_2043:item
  food_bacon_2044:item
  food_banana_2045:item
  food_cake_2046:item
  food_carrot_2047:item
  food_cereal_2048:item
  food_cheese_2049:item
  food_chicken_2050:item
  food_dessert_2051:item
  food_donut_2052:item
  food_egg_2053:item
  food_fish_2054:item
  food_food_2055:item
  food_fruit_2056:item
  food_hamburger_2057:item
  food_ice_cream_2058:item
  food_jam_2059:item
  food_kiwi_2060:item
  food_lemon_2061:item
  food_noodles_2062:item
  food_oatmeal_2063:item
  food_peanut_butter_2064:item
  food_pizza_2065:item
  food_potato_2066:item
  food_rice_2067:item
  food_salt_2068:item
  food_snack_2069:item
  food_sugar_2070:item
  food_turkey_2071:item
  food_vegetable_2072:item
  dry_pasta_2073:item
  milk_2074:item
  clothes_dress_2075:item
  clothes_hat_2076:item
  clothes_gloves_2077:item
  clothes_jacket_2078:item
  clothes_scarf_2079:item
  cutting_board_2080:item
  remote_control_2081:item
  cat_2082:item
  towel_2083:item
  cd_player_2084:item
  dvd_player_2085:item
  headset_2086:item
  cup_2087:item
  cup_2088:item
  cup_2089:item
  stove_2090:item
  book_2091:item
  book_2092:item
  pot_2093:item
  vacuum_cleaner_2094:item
  bowl_2095:item
  bowl_2096:item
  bowl_2097:item
  cleaning_solution_2098:item
  ironing_board_2099:item
  cd_2100:item
  sauce_2101:item
  oil_2102:item
  fork_2103:item
  fork_2104:item
  plate_2105:item
  spectacles_2106:item
  fryingpan_2107:item
  detergent_2108:item
  window_2109:item
  computer_2110:item
  dining_room_1:item
  wall_2:item
  wall_3:item
  wall_4:item
  wall_5:item
  wall_6:item
  wall_7:item
  wall_8:item
  wall_9:item
  wall_10:item
  wall_11:item
  floor_12:item
  floor_13:item
  floor_14:item
  floor_15:item
  floor_16:item
  floor_17:item
  floor_18:item
  floor_19:item
  floor_20:item
  floor_21:item
  floor_22:item
  floor_23:item
  floor_24:item
  ceiling_25:item
  ceiling_26:item
  ceiling_27:item
  ceiling_28:item
  ceiling_29:item
  ceiling_30:item
  ceiling_31:item
  ceiling_32:item
  ceiling_33:item
  ceiling_34:item
  ceiling_35:item
  ceiling_36:item
  doorjamb_37:item
  door_38:item
  doorjamb_39:item
  window_40:item
  ceilinglamp_41:item
  ceilinglamp_42:item
  ceilinglamp_43:item
  walllamp_44:item
  walllamp_45:item
  walllamp_46:item
  phone_47:item
  powersocket_48:item
  light_49:item
  knifeblock_52:item
  pot_54:item
  photoframe_102:item
  mat_114:item
  mat_115:item
  orchid_117:item
  drawing_118:item
  curtain_119:item
  curtain_120:item
  curtain_121:item
  bench_122:item
  table_123:item
  bench_124:item
  bench_125:item
  bench_126:item
  table_127:item
  kitchen_counter_128:item
  kitchen_counter_129:item
  cupboard_130:item
  cupboard_131:item
  kitchen_counter_132:item
  sink_133:item
  faucet_134:item
  tvstand_135:item
  bookshelf_136:item
  bookshelf_137:item
  chair_138:item
  stovefan_139:item
  fridge_140:item
  oven_141:item
  tray_142:item
  dishwasher_143:item
  toaster_144:item
  coffe_maker_147:item
  microwave_149:item
  home_office_161:item
  floor_162:item
  floor_163:item
  floor_164:item
  floor_165:item
  floor_166:item
  floor_167:item
  floor_168:item
  wall_169:item
  wall_170:item
  wall_171:item
  wall_172:item
  wall_173:item
  wall_174:item
  ceiling_175:item
  ceiling_176:item
  ceiling_177:item
  ceiling_178:item
  ceiling_179:item
  ceiling_180:item
  window_181:item
  doorjamb_182:item
  walllamp_183:item
  walllamp_184:item
  ceilinglamp_185:item
  tvstand_186:item
  wallshelf_187:item
  bookshelf_188:item
  bookshelf_189:item
  wallshelf_190:item
  wallshelf_191:item
  couch_192:item
  table_193:item
  pillow_195:item
  drawing_196:item
  curtain_197:item
  curtain_198:item
  curtain_199:item
  orchid_200:item
  mat_201:item
  photoframe_210:item
  television_216:item
  light_217:item
  powersocket_218:item
  bedroom_220:item
  floor_221:item
  floor_222:item
  floor_223:item
  floor_224:item
  floor_225:item
  ceiling_226:item
  ceiling_227:item
  ceiling_228:item
  ceiling_229:item
  wall_230:item
  wall_231:item
  wall_232:item
  wall_233:item
  door_234:item
  ceilinglamp_235:item
  tablelamp_236:item
  mat_237:item
  drawing_238:item
  pillow_239:item
  pillow_240:item
  photoframe_246:item
  light_258:item
  powersocket_259:item
  bookshelf_260:item
  desk_261:item
  nightstand_262:item
  chair_263:item
  bed_264:item
  bathroom_265:item
  wall_266:item
  wall_267:item
  wall_268:item
  wall_269:item
  wall_270:item
  wall_271:item
  floor_272:item
  floor_273:item
  floor_274:item
  floor_275:item
  floor_276:item
  floor_277:item
  floor_278:item
  ceiling_279:item
  ceiling_280:item
  ceiling_281:item
  ceiling_282:item
  ceiling_283:item
  ceiling_284:item
  doorjamb_285:item
  door_286:item
  window_287:item
  ceilinglamp_288:item
  walllamp_289:item
  walllamp_290:item
  walllamp_291:item
  mat_292:item
  curtain_293:item
  curtain_294:item
  drawing_296:item
  bathtub_297:item
  towel_rack_298:item
  towel_rack_299:item
  towel_rack_300:item
  wallshelf_301:item
  toilet_302:item
  shower_303:item
  curtain_304:item
  bathroom_cabinet_305:item
  bathroom_counter_306:item
  sink_307:item
  faucet_308:item
  light_325:item
  bedroom_327:item
  floor_328:item
  floor_329:item
  floor_330:item
  floor_331:item
  floor_332:item
  floor_333:item
  floor_334:item
  floor_335:item
  floor_336:item
  floor_337:item
  wall_338:item
  wall_339:item
  wall_340:item
  wall_341:item
  wall_342:item
  wall_343:item
  wall_344:item
  wall_345:item
  window_346:item
  ceiling_347:item
  ceiling_348:item
  ceiling_349:item
  ceiling_350:item
  ceiling_351:item
  ceiling_352:item
  ceiling_353:item
  ceiling_354:item
  ceiling_355:item
  doorjamb_356:item
  ceilinglamp_357:item
  tablelamp_358:item
  tablelamp_359:item
  trashcan_360:item
  photoframe_361:item
  pillow_368:item
  pillow_370:item
  bookshelf_372:item
  nightstand_373:item
  chair_374:item
  desk_375:item
  bed_376:item
  dresser_377:item
  filing_cabinet_378:item
  computer_379:item
  mouse_380:item
  mousepad_381:item
  keyboard_382:item
  cpuscreen_383:item
  light_384:item
  mat_386:item
  drawing_387:item
  drawing_388:item
  drawing_389:item
  curtain_390:item
  curtain_391:item
  curtain_392:item
  dvd_player_2000:item
  shoes_2001:item
  alcohol_2002:item
  mouse_2003:item
  coin_2004:item
  oil_2005:item
  cup_2006:item
  stereo_2007:item
  food_orange_2008:item
  bills_2009:item
  novel_2010:item
  homework_2011:item
  needle_2012:item
  glue_2013:item
  napkin_2014:item
  laptop_2015:item
  food_bread_2016:item
  tea_bag_2017:item
  food_butter_2018:item
  video_game_controller_2019:item
  crayon_2020:item
  dough_2021:item
  clothes_underwear_2022:item
  box_2023:item
  needle_2024:item
  laser_pointer_2025:item
  food_onion_2026:item
  console_2027:item
  tape_2028:item
  after_shave_2029:item
  crayon_2030:item
  stamp_2031:item
  blender_2032:item
  check_2033:item
  juice_2034:item
  coffee_filter_2035:item
  knife_2036:item
  soap_2037:item
  soap_2038:item
  pajamas_2039:item
#object_end

init:
    #categories
    is_keyboard[keyboard_2111]=True
    is_mouse[mouse_2112]=True
    is_clothes_pants[clothes_pants_2113]=True
    is_pants[clothes_pants_2113]=True
    is_clothes_shirt[clothes_shirt_2114]=True
    is_shirt[clothes_shirt_2114]=True
    is_clothes_socks[clothes_socks_2115]=True
    is_clothes_skirt[clothes_skirt_2116]=True
    is_iron[iron_2117]=True
    is_chair[chair_2118]=True
    is_basket_for_clothes[basket_for_clothes_2040]=True
    is_clothes_pile[basket_for_clothes_2040]=True
    is_washing_machine[washing_machine_2041]=True
    is_food_steak[food_steak_2042]=True
    is_apple[food_apple_2043]=True
    is_food_apple[food_apple_2043]=True
    is_food_bacon[food_bacon_2044]=True
    is_banana[food_banana_2045]=True
    is_food_banana[food_banana_2045]=True
    is_food_cake[food_cake_2046]=True
    is_food_carrot[food_carrot_2047]=True
    is_carrot[food_carrot_2047]=True
    is_food_cereal[food_cereal_2048]=True
    is_cereal[food_cereal_2048]=True
    is_food_cheese[food_cheese_2049]=True
    is_chicken[food_chicken_2050]=True
    is_food_chicken[food_chicken_2050]=True
    is_poundcake[food_dessert_2051]=True
    is_pie[food_dessert_2051]=True
    is_pudding[food_dessert_2051]=True
    is_pancake[food_dessert_2051]=True
    is_milkshake[food_dessert_2051]=True
    is_watermelon[food_dessert_2051]=True
    is_cupcake[food_dessert_2051]=True
    is_creamybuns[food_dessert_2051]=True
    is_sundae[food_dessert_2051]=True
    is_food_dessert[food_dessert_2051]=True
    is_food_donut[food_donut_2052]=True
    is_food_egg[food_egg_2053]=True
    is_salmon[food_fish_2054]=True
    is_food_fish[food_fish_2054]=True
    is_bellpepper[food_food_2055]=True
    is_apple[food_food_2055]=True
    is_tomato[food_food_2055]=True
    is_cutlets[food_food_2055]=True
    is_whippedcream[food_food_2055]=True
    is_crackers[food_food_2055]=True
    is_potato[food_food_2055]=True
    is_plum[food_food_2055]=True
    is_banana[food_food_2055]=True
    is_bananas[food_food_2055]=True
    is_food_food[food_food_2055]=True
    is_creamybuns[food_food_2055]=True
    is_chicken[food_food_2055]=True
    is_pear[food_food_2055]=True
    is_cereal[food_food_2055]=True
    is_salmon[food_food_2055]=True
    is_bell_pepper[food_food_2055]=True
    is_chocolatesyrup[food_food_2055]=True
    is_chinesefood[food_food_2055]=True
    is_orange[food_food_2055]=True
    is_cucumber[food_food_2055]=True
    is_pear[food_fruit_2056]=True
    is_apple[food_fruit_2056]=True
    is_plum[food_fruit_2056]=True
    is_banana[food_fruit_2056]=True
    is_orange[food_fruit_2056]=True
    is_food_fruit[food_fruit_2056]=True
    is_watermelon[food_fruit_2056]=True
    is_mincedmeat[food_hamburger_2057]=True
    is_food_hamburger[food_hamburger_2057]=True
    is_food_ice_cream[food_ice_cream_2058]=True
    is_food_jam[food_jam_2059]=True
    is_food_kiwi[food_kiwi_2060]=True
    is_lemon[food_lemon_2061]=True
    is_food_lemon[food_lemon_2061]=True
    is_food_noodles[food_noodles_2062]=True
    is_food_oatmeal[food_oatmeal_2063]=True
    is_cereal[food_oatmeal_2063]=True
    is_food_peanut_butter[food_peanut_butter_2064]=True
    is_food_pizza[food_pizza_2065]=True
    is_food_potato[food_potato_2066]=True
    is_potato[food_potato_2066]=True
    is_food_rice[food_rice_2067]=True
    is_food_salt[food_salt_2068]=True
    is_condiment_shaker[food_salt_2068]=True
    is_poundcake[food_snack_2069]=True
    is_chips[food_snack_2069]=True
    is_food_snack[food_snack_2069]=True
    is_crackers[food_snack_2069]=True
    is_apple[food_snack_2069]=True
    is_salt_crackers[food_snack_2069]=True
    is_candybar[food_snack_2069]=True
    is_banana[food_snack_2069]=True
    is_cupcake[food_snack_2069]=True
    is_food_sugar[food_sugar_2070]=True
    is_condiment_shaker[food_sugar_2070]=True
    is_food_turkey[food_turkey_2071]=True
    is_chicken[food_turkey_2071]=True
    is_salad[food_vegetable_2072]=True
    is_carrot[food_vegetable_2072]=True
    is_tomato[food_vegetable_2072]=True
    is_potato[food_vegetable_2072]=True
    is_food_vegetable[food_vegetable_2072]=True
    is_cucumber[food_vegetable_2072]=True
    is_dry_pasta[dry_pasta_2073]=True
    is_milk[milk_2074]=True
    is_clothes_dress[clothes_dress_2075]=True
    is_clothes_hat[clothes_hat_2076]=True
    is_clothes_gloves[clothes_gloves_2077]=True
    is_clothes_jacket[clothes_jacket_2078]=True
    is_clothes_scarf[clothes_scarf_2079]=True
    is_cutting_board[cutting_board_2080]=True
    is_controller[remote_control_2081]=True
    is_remote_control[remote_control_2081]=True
    is_cat[cat_2082]=True
    is_towel[towel_2083]=True
    is_radio[cd_player_2084]=True
    is_cd_player[cd_player_2084]=True
    is_dvd_player[dvd_player_2085]=True
    is_headset[headset_2086]=True
    is_cup[cup_2087]=True
    is_mug[cup_2087]=True
    is_wineglass[cup_2087]=True
    is_waterglass[cup_2087]=True
    is_cup[cup_2088]=True
    is_mug[cup_2088]=True
    is_wineglass[cup_2088]=True
    is_waterglass[cup_2088]=True
    is_cup[cup_2089]=True
    is_mug[cup_2089]=True
    is_wineglass[cup_2089]=True
    is_waterglass[cup_2089]=True
    is_stove[stove_2090]=True
    is_oven[stove_2090]=True
    is_textbook[book_2091]=True
    is_book[book_2091]=True
    is_novel[book_2091]=True
    is_textbook[book_2092]=True
    is_book[book_2092]=True
    is_novel[book_2092]=True
    is_pot[pot_2093]=True
    is_vacuum_cleaner[vacuum_cleaner_2094]=True
    is_bowl[bowl_2095]=True
    is_dish_bowl[bowl_2095]=True
    is_bowl[bowl_2096]=True
    is_dish_bowl[bowl_2096]=True
    is_bowl[bowl_2097]=True
    is_dish_bowl[bowl_2097]=True
    is_dishwashingliquid[cleaning_solution_2098]=True
    is_cleaning_solution[cleaning_solution_2098]=True
    is_ironing_board[ironing_board_2099]=True
    is_cd[cd_2100]=True
    is_sauce[sauce_2101]=True
    is_condiment_bottle[sauce_2101]=True
    is_oil[oil_2102]=True
    is_condiment_bottle[oil_2102]=True
    is_fork[fork_2103]=True
    is_cutlery_fork[fork_2103]=True
    is_fork[fork_2104]=True
    is_cutlery_fork[fork_2104]=True
    is_plate[plate_2105]=True
    is_glasses[spectacles_2106]=True
    is_spectacles[spectacles_2106]=True
    is_fryingpan[fryingpan_2107]=True
    is_detergent[detergent_2108]=True
    is_dishwashingliquid[detergent_2108]=True
    is_window[window_2109]=True
    is_pc[computer_2110]=True
    is_cpu_case[computer_2110]=True
    is_computer[computer_2110]=True
    is_dining_room[dining_room_1]=True
    is_kitchen[dining_room_1]=True
    is_wall[wall_2]=True
    is_wall[wall_3]=True
    is_wall[wall_4]=True
    is_wall[wall_5]=True
    is_wall[wall_6]=True
    is_wall[wall_7]=True
    is_wall[wall_8]=True
    is_wall[wall_9]=True
    is_wall[wall_10]=True
    is_wall[wall_11]=True
    is_floor[floor_12]=True
    is_floor[floor_13]=True
    is_floor[floor_14]=True
    is_floor[floor_15]=True
    is_floor[floor_16]=True
    is_floor[floor_17]=True
    is_floor[floor_18]=True
    is_floor[floor_19]=True
    is_floor[floor_20]=True
    is_floor[floor_21]=True
    is_floor[floor_22]=True
    is_floor[floor_23]=True
    is_floor[floor_24]=True
    is_ceiling[ceiling_25]=True
    is_ceiling[ceiling_26]=True
    is_ceiling[ceiling_27]=True
    is_ceiling[ceiling_28]=True
    is_ceiling[ceiling_29]=True
    is_ceiling[ceiling_30]=True
    is_ceiling[ceiling_31]=True
    is_ceiling[ceiling_32]=True
    is_ceiling[ceiling_33]=True
    is_ceiling[ceiling_34]=True
    is_ceiling[ceiling_35]=True
    is_ceiling[ceiling_36]=True
    is_doorjamb[doorjamb_37]=True
    is_door[door_38]=True
    is_doorjamb[doorjamb_39]=True
    is_window[window_40]=True
    is_ceilinglamp[ceilinglamp_41]=True
    is_ceilinglamp[ceilinglamp_42]=True
    is_ceilinglamp[ceilinglamp_43]=True
    is_walllamp[walllamp_44]=True
    is_walllamp[walllamp_45]=True
    is_walllamp[walllamp_46]=True
    is_cellphone[phone_47]=True
    is_wall_phone[phone_47]=True
    is_phone[phone_47]=True
    is_powersocket[powersocket_48]=True
    is_light[light_49]=True
    is_light_switch[light_49]=True
    is_lightswitch[light_49]=True
    is_knifeblock[knifeblock_52]=True
    is_pot[pot_54]=True
    is_photoframe[photoframe_102]=True
    is_rug[mat_114]=True
    is_mat[mat_114]=True
    is_rug[mat_115]=True
    is_mat[mat_115]=True
    is_orchid[orchid_117]=True
    is_drawing[drawing_118]=True
    is_wallpictureframe[drawing_118]=True
    is_curtain[curtain_119]=True
    is_curtains[curtain_119]=True
    is_curtain[curtain_120]=True
    is_curtains[curtain_120]=True
    is_curtain[curtain_121]=True
    is_curtains[curtain_121]=True
    is_bench[bench_122]=True
    is_table[table_123]=True
    is_diningtable[table_123]=True
    is_coffee_table[table_123]=True
    is_kitchen_table[table_123]=True
    is_bench[bench_124]=True
    is_bench[bench_125]=True
    is_bench[bench_126]=True
    is_table[table_127]=True
    is_diningtable[table_127]=True
    is_coffee_table[table_127]=True
    is_kitchen_table[table_127]=True
    is_kitchen_counter[kitchen_counter_128]=True
    is_kitchen_counter[kitchen_counter_129]=True
    is_kitchen_cabinets[cupboard_130]=True
    is_cupboard[cupboard_130]=True
    is_kitchen_cabinets[cupboard_131]=True
    is_cupboard[cupboard_131]=True
    is_kitchen_counter[kitchen_counter_132]=True
    is_sink[sink_133]=True
    is_faucet[faucet_134]=True
    is_tvstand[tvstand_135]=True
    is_bookshelf[bookshelf_136]=True
    is_bookshelf[bookshelf_137]=True
    is_chair[chair_138]=True
    is_stovefan[stovefan_139]=True
    is_freezer[fridge_140]=True
    is_fridge[fridge_140]=True
    is_stove[oven_141]=True
    is_oven[oven_141]=True
    is_oventray[tray_142]=True
    is_tray[tray_142]=True
    is_dishwasher[dishwasher_143]=True
    is_toaster[toaster_144]=True
    is_coffe_maker[coffe_maker_147]=True
    is_coffeemaker[coffe_maker_147]=True
    is_microwave[microwave_149]=True
    is_home_office[home_office_161]=True
    is_livingroom[home_office_161]=True
    is_floor[floor_162]=True
    is_floor[floor_163]=True
    is_floor[floor_164]=True
    is_floor[floor_165]=True
    is_floor[floor_166]=True
    is_floor[floor_167]=True
    is_floor[floor_168]=True
    is_wall[wall_169]=True
    is_wall[wall_170]=True
    is_wall[wall_171]=True
    is_wall[wall_172]=True
    is_wall[wall_173]=True
    is_wall[wall_174]=True
    is_ceiling[ceiling_175]=True
    is_ceiling[ceiling_176]=True
    is_ceiling[ceiling_177]=True
    is_ceiling[ceiling_178]=True
    is_ceiling[ceiling_179]=True
    is_ceiling[ceiling_180]=True
    is_window[window_181]=True
    is_doorjamb[doorjamb_182]=True
    is_walllamp[walllamp_183]=True
    is_walllamp[walllamp_184]=True
    is_ceilinglamp[ceilinglamp_185]=True
    is_tvstand[tvstand_186]=True
    is_wallshelf[wallshelf_187]=True
    is_bookshelf[bookshelf_188]=True
    is_bookshelf[bookshelf_189]=True
    is_wallshelf[wallshelf_190]=True
    is_wallshelf[wallshelf_191]=True
    is_couch[couch_192]=True
    is_sofa[couch_192]=True
    is_table[table_193]=True
    is_diningtable[table_193]=True
    is_coffee_table[table_193]=True
    is_kitchen_table[table_193]=True
    is_pillow[pillow_195]=True
    is_drawing[drawing_196]=True
    is_wallpictureframe[drawing_196]=True
    is_curtain[curtain_197]=True
    is_curtains[curtain_197]=True
    is_curtain[curtain_198]=True
    is_curtains[curtain_198]=True
    is_curtain[curtain_199]=True
    is_curtains[curtain_199]=True
    is_orchid[orchid_200]=True
    is_rug[mat_201]=True
    is_mat[mat_201]=True
    is_photoframe[photoframe_210]=True
    is_tv[television_216]=True
    is_walltv[television_216]=True
    is_television[television_216]=True
    is_light[light_217]=True
    is_light_switch[light_217]=True
    is_lightswitch[light_217]=True
    is_powersocket[powersocket_218]=True
    is_bedroom[bedroom_220]=True
    is_floor[floor_221]=True
    is_floor[floor_222]=True
    is_floor[floor_223]=True
    is_floor[floor_224]=True
    is_floor[floor_225]=True
    is_ceiling[ceiling_226]=True
    is_ceiling[ceiling_227]=True
    is_ceiling[ceiling_228]=True
    is_ceiling[ceiling_229]=True
    is_wall[wall_230]=True
    is_wall[wall_231]=True
    is_wall[wall_232]=True
    is_wall[wall_233]=True
    is_door[door_234]=True
    is_ceilinglamp[ceilinglamp_235]=True
    is_tablelamp[tablelamp_236]=True
    is_rug[mat_237]=True
    is_mat[mat_237]=True
    is_drawing[drawing_238]=True
    is_wallpictureframe[drawing_238]=True
    is_pillow[pillow_239]=True
    is_pillow[pillow_240]=True
    is_photoframe[photoframe_246]=True
    is_light[light_258]=True
    is_light_switch[light_258]=True
    is_lightswitch[light_258]=True
    is_powersocket[powersocket_259]=True
    is_bookshelf[bookshelf_260]=True
    is_cpu_table[desk_261]=True
    is_desk[desk_261]=True
    is_nightstand[nightstand_262]=True
    is_chair[chair_263]=True
    is_bed[bed_264]=True
    is_bathroom[bathroom_265]=True
    is_wall[wall_266]=True
    is_wall[wall_267]=True
    is_wall[wall_268]=True
    is_wall[wall_269]=True
    is_wall[wall_270]=True
    is_wall[wall_271]=True
    is_floor[floor_272]=True
    is_floor[floor_273]=True
    is_floor[floor_274]=True
    is_floor[floor_275]=True
    is_floor[floor_276]=True
    is_floor[floor_277]=True
    is_floor[floor_278]=True
    is_ceiling[ceiling_279]=True
    is_ceiling[ceiling_280]=True
    is_ceiling[ceiling_281]=True
    is_ceiling[ceiling_282]=True
    is_ceiling[ceiling_283]=True
    is_ceiling[ceiling_284]=True
    is_doorjamb[doorjamb_285]=True
    is_door[door_286]=True
    is_window[window_287]=True
    is_ceilinglamp[ceilinglamp_288]=True
    is_walllamp[walllamp_289]=True
    is_walllamp[walllamp_290]=True
    is_walllamp[walllamp_291]=True
    is_rug[mat_292]=True
    is_mat[mat_292]=True
    is_curtain[curtain_293]=True
    is_curtains[curtain_293]=True
    is_curtain[curtain_294]=True
    is_curtains[curtain_294]=True
    is_drawing[drawing_296]=True
    is_wallpictureframe[drawing_296]=True
    is_bathtub[bathtub_297]=True
    is_towel_rack[towel_rack_298]=True
    is_towel_rack[towel_rack_299]=True
    is_towel_rack[towel_rack_300]=True
    is_wallshelf[wallshelf_301]=True
    is_toilet[toilet_302]=True
    is_shower[shower_303]=True
    is_stall[shower_303]=True
    is_curtain[curtain_304]=True
    is_curtains[curtain_304]=True
    is_bathroom_cabinet[bathroom_cabinet_305]=True
    is_bathroom_counter[bathroom_counter_306]=True
    is_sink[sink_307]=True
    is_faucet[faucet_308]=True
    is_light[light_325]=True
    is_light_switch[light_325]=True
    is_lightswitch[light_325]=True
    is_bedroom[bedroom_327]=True
    is_floor[floor_328]=True
    is_floor[floor_329]=True
    is_floor[floor_330]=True
    is_floor[floor_331]=True
    is_floor[floor_332]=True
    is_floor[floor_333]=True
    is_floor[floor_334]=True
    is_floor[floor_335]=True
    is_floor[floor_336]=True
    is_floor[floor_337]=True
    is_wall[wall_338]=True
    is_wall[wall_339]=True
    is_wall[wall_340]=True
    is_wall[wall_341]=True
    is_wall[wall_342]=True
    is_wall[wall_343]=True
    is_wall[wall_344]=True
    is_wall[wall_345]=True
    is_window[window_346]=True
    is_ceiling[ceiling_347]=True
    is_ceiling[ceiling_348]=True
    is_ceiling[ceiling_349]=True
    is_ceiling[ceiling_350]=True
    is_ceiling[ceiling_351]=True
    is_ceiling[ceiling_352]=True
    is_ceiling[ceiling_353]=True
    is_ceiling[ceiling_354]=True
    is_ceiling[ceiling_355]=True
    is_doorjamb[doorjamb_356]=True
    is_ceilinglamp[ceilinglamp_357]=True
    is_tablelamp[tablelamp_358]=True
    is_tablelamp[tablelamp_359]=True
    is_trashcan[trashcan_360]=True
    is_garbage_can[trashcan_360]=True
    is_photoframe[photoframe_361]=True
    is_pillow[pillow_368]=True
    is_pillow[pillow_370]=True
    is_bookshelf[bookshelf_372]=True
    is_nightstand[nightstand_373]=True
    is_chair[chair_374]=True
    is_cpu_table[desk_375]=True
    is_desk[desk_375]=True
    is_bed[bed_376]=True
    is_closet[dresser_377]=True
    is_dresser[dresser_377]=True
    is_cabinet[filing_cabinet_378]=True
    is_filing_cabinet[filing_cabinet_378]=True
    is_pc[computer_379]=True
    is_cpu_case[computer_379]=True
    is_computer[computer_379]=True
    is_mouse[mouse_380]=True
    is_mousemat[mousepad_381]=True
    is_mouse_mat[mousepad_381]=True
    is_mousepad[mousepad_381]=True
    is_keyboard[keyboard_382]=True
    is_cpuscreen[cpuscreen_383]=True
    is_light[light_384]=True
    is_light_switch[light_384]=True
    is_lightswitch[light_384]=True
    is_rug[mat_386]=True
    is_mat[mat_386]=True
    is_drawing[drawing_387]=True
    is_wallpictureframe[drawing_387]=True
    is_drawing[drawing_388]=True
    is_wallpictureframe[drawing_388]=True
    is_drawing[drawing_389]=True
    is_wallpictureframe[drawing_389]=True
    is_curtain[curtain_390]=True
    is_curtains[curtain_390]=True
    is_curtain[curtain_391]=True
    is_curtains[curtain_391]=True
    is_curtain[curtain_392]=True
    is_curtains[curtain_392]=True
    is_dvd_player[dvd_player_2000]=True
    is_shoes[shoes_2001]=True
    is_slippers[shoes_2001]=True
    is_alcohol[alcohol_2002]=True
    is_mouse[mouse_2003]=True
    is_coin[coin_2004]=True
    is_oil[oil_2005]=True
    is_condiment_bottle[oil_2005]=True
    is_cup[cup_2006]=True
    is_mug[cup_2006]=True
    is_wineglass[cup_2006]=True
    is_waterglass[cup_2006]=True
    is_radio[stereo_2007]=True
    is_stereo[stereo_2007]=True
    is_food_orange[food_orange_2008]=True
    is_bills[bills_2009]=True
    is_book[novel_2010]=True
    is_novel[novel_2010]=True
    is_homework[homework_2011]=True
    is_needle[needle_2012]=True
    is_glue[glue_2013]=True
    is_papertowel[napkin_2014]=True
    is_cloth_napkin[napkin_2014]=True
    is_napkin[napkin_2014]=True
    is_laptop[laptop_2015]=True
    is_food_bread[food_bread_2016]=True
    is_bread_slice[food_bread_2016]=True
    is_bread[food_bread_2016]=True
    is_tea_bag[tea_bag_2017]=True
    is_food_butter[food_butter_2018]=True
    is_video_game_controller[video_game_controller_2019]=True
    is_crayon[crayon_2020]=True
    is_crayons[crayon_2020]=True
    is_dough[dough_2021]=True
    is_clothes_underwear[clothes_underwear_2022]=True
    is_box[box_2023]=True
    is_needle[needle_2024]=True
    is_laser_pointer[laser_pointer_2025]=True
    is_food_onion[food_onion_2026]=True
    is_console[console_2027]=True
    is_tape[tape_2028]=True
    is_face_cream[after_shave_2029]=True
    is_after_shave[after_shave_2029]=True
    is_facecream[after_shave_2029]=True
    is_crayon[crayon_2030]=True
    is_crayons[crayon_2030]=True
    is_stamp[stamp_2031]=True
    is_blender[blender_2032]=True
    is_check[check_2033]=True
    is_paper[check_2033]=True
    is_juice[juice_2034]=True
    is_coffee_filter[coffee_filter_2035]=True
    is_chefknife[knife_2036]=True
    is_cutlery_knife[knife_2036]=True
    is_knife[knife_2036]=True
    is_barsoap[soap_2037]=True
    is_soap[soap_2037]=True
    is_barsoap[soap_2038]=True
    is_soap[soap_2038]=True
    is_pajamas[pajamas_2039]=True
    #categories_end

    #states
    is_on[ceilinglamp_41]=True
    is_on[ceilinglamp_42]=True
    is_on[ceilinglamp_43]=True
    is_on[walllamp_44]=True
    is_on[walllamp_45]=True
    is_on[walllamp_46]=True
    is_on[faucet_134]=True
    is_on[fridge_140]=True
    is_on[walllamp_183]=True
    is_on[walllamp_184]=True
    is_on[ceilinglamp_185]=True
    is_on[ceilinglamp_235]=True
    is_on[tablelamp_236]=True
    is_on[ceilinglamp_288]=True
    is_on[walllamp_289]=True
    is_on[walllamp_290]=True
    is_on[walllamp_291]=True
    is_on[faucet_308]=True
    is_on[ceilinglamp_357]=True
    is_on[tablelamp_358]=True
    is_on[tablelamp_359]=True
    is_off[washing_machine_2041]=True
    is_off[stove_2090]=True
    is_off[computer_2110]=True
    is_off[light_49]=True
    is_off[oven_141]=True
    is_off[dishwasher_143]=True
    is_off[toaster_144]=True
    is_off[coffe_maker_147]=True
    is_off[microwave_149]=True
    is_off[television_216]=True
    is_off[light_217]=True
    is_off[light_258]=True
    is_off[toilet_302]=True
    is_off[shower_303]=True
    is_off[light_325]=True
    is_off[computer_379]=True
    is_off[light_384]=True
    open[doorjamb_37]=True
    open[door_38]=True
    open[doorjamb_39]=True
    open[cupboard_130]=True
    open[kitchen_counter_132]=True
    open[bookshelf_136]=True
    open[doorjamb_182]=True
    open[door_234]=True
    open[nightstand_262]=True
    open[doorjamb_285]=True
    open[door_286]=True
    open[doorjamb_356]=True
    open[trashcan_360]=True
    open[nightstand_373]=True
    open[dresser_377]=True
    open[filing_cabinet_378]=True
    open[curtain_391]=True
    closed[washing_machine_2041]=True
    closed[stove_2090]=True
    closed[window_2109]=True
    closed[window_40]=True
    closed[light_49]=True
    closed[curtain_119]=True
    closed[curtain_120]=True
    closed[curtain_121]=True
    closed[kitchen_counter_128]=True
    closed[kitchen_counter_129]=True
    closed[cupboard_131]=True
    closed[bookshelf_137]=True
    closed[fridge_140]=True
    closed[oven_141]=True
    closed[dishwasher_143]=True
    closed[coffe_maker_147]=True
    closed[microwave_149]=True
    closed[window_181]=True
    closed[bookshelf_188]=True
    closed[bookshelf_189]=True
    closed[curtain_197]=True
    closed[curtain_198]=True
    closed[curtain_199]=True
    closed[light_217]=True
    closed[light_258]=True
    closed[bookshelf_260]=True
    closed[window_287]=True
    closed[curtain_293]=True
    closed[curtain_294]=True
    closed[toilet_302]=True
    closed[curtain_304]=True
    closed[bathroom_cabinet_305]=True
    closed[bathroom_counter_306]=True
    closed[light_325]=True
    closed[window_346]=True
    closed[bookshelf_372]=True
    closed[light_384]=True
    closed[curtain_390]=True
    closed[curtain_392]=True
    dirty[window_2109]=True
    dirty[wall_2]=True
    dirty[wall_3]=True
    dirty[wall_4]=True
    dirty[wall_8]=True
    dirty[wall_9]=True
    dirty[wall_11]=True
    dirty[floor_12]=True
    dirty[floor_13]=True
    dirty[floor_17]=True
    dirty[floor_18]=True
    dirty[floor_21]=True
    dirty[floor_22]=True
    dirty[floor_24]=True
    dirty[ceiling_26]=True
    dirty[ceiling_27]=True
    dirty[ceiling_29]=True
    dirty[ceiling_30]=True
    dirty[ceiling_31]=True
    dirty[ceiling_35]=True
    dirty[ceiling_36]=True
    dirty[window_40]=True
    dirty[sink_133]=True
    dirty[floor_164]=True
    dirty[floor_165]=True
    dirty[floor_168]=True
    dirty[wall_170]=True
    dirty[wall_171]=True
    dirty[ceiling_175]=True
    dirty[ceiling_176]=True
    dirty[window_181]=True
    dirty[bookshelf_188]=True
    dirty[floor_221]=True
    dirty[floor_225]=True
    dirty[ceiling_227]=True
    dirty[ceiling_228]=True
    dirty[wall_233]=True
    dirty[wall_266]=True
    dirty[wall_270]=True
    dirty[floor_273]=True
    dirty[floor_276]=True
    dirty[floor_277]=True
    dirty[floor_278]=True
    dirty[ceiling_281]=True
    dirty[ceiling_282]=True
    dirty[ceiling_283]=True
    dirty[window_287]=True
    dirty[curtain_293]=True
    dirty[curtain_294]=True
    dirty[bathroom_cabinet_305]=True
    dirty[sink_307]=True
    dirty[floor_328]=True
    dirty[floor_329]=True
    dirty[floor_331]=True
    dirty[floor_332]=True
    dirty[floor_333]=True
    dirty[floor_335]=True
    dirty[wall_338]=True
    dirty[wall_339]=True
    dirty[window_346]=True
    dirty[ceiling_350]=True
    dirty[ceiling_352]=True
    dirty[ceiling_353]=True
    clean[washing_machine_2041]=True
    clean[cutting_board_2080]=True
    clean[computer_2110]=True
    clean[dining_room_1]=True
    clean[wall_5]=True
    clean[wall_6]=True
    clean[wall_7]=True
    clean[wall_10]=True
    clean[floor_14]=True
    clean[floor_15]=True
    clean[floor_16]=True
    clean[floor_19]=True
    clean[floor_20]=True
    clean[floor_23]=True
    clean[ceiling_25]=True
    clean[ceiling_28]=True
    clean[ceiling_32]=True
    clean[ceiling_33]=True
    clean[ceiling_34]=True
    clean[doorjamb_37]=True
    clean[door_38]=True
    clean[doorjamb_39]=True
    clean[ceilinglamp_41]=True
    clean[ceilinglamp_42]=True
    clean[ceilinglamp_43]=True
    clean[walllamp_44]=True
    clean[walllamp_45]=True
    clean[walllamp_46]=True
    clean[powersocket_48]=True
    clean[light_49]=True
    clean[knifeblock_52]=True
    clean[photoframe_102]=True
    clean[orchid_117]=True
    clean[curtain_119]=True
    clean[curtain_120]=True
    clean[curtain_121]=True
    clean[bench_122]=True
    clean[table_123]=True
    clean[bench_124]=True
    clean[bench_125]=True
    clean[bench_126]=True
    clean[table_127]=True
    clean[kitchen_counter_128]=True
    clean[kitchen_counter_129]=True
    clean[cupboard_130]=True
    clean[cupboard_131]=True
    clean[kitchen_counter_132]=True
    clean[faucet_134]=True
    clean[tvstand_135]=True
    clean[bookshelf_136]=True
    clean[bookshelf_137]=True
    clean[stovefan_139]=True
    clean[fridge_140]=True
    clean[oven_141]=True
    clean[dishwasher_143]=True
    clean[toaster_144]=True
    clean[coffe_maker_147]=True
    clean[microwave_149]=True
    clean[home_office_161]=True
    clean[floor_162]=True
    clean[floor_163]=True
    clean[floor_166]=True
    clean[floor_167]=True
    clean[wall_169]=True
    clean[wall_172]=True
    clean[wall_173]=True
    clean[wall_174]=True
    clean[ceiling_177]=True
    clean[ceiling_178]=True
    clean[ceiling_179]=True
    clean[ceiling_180]=True
    clean[doorjamb_182]=True
    clean[walllamp_183]=True
    clean[walllamp_184]=True
    clean[ceilinglamp_185]=True
    clean[tvstand_186]=True
    clean[wallshelf_187]=True
    clean[bookshelf_189]=True
    clean[wallshelf_190]=True
    clean[wallshelf_191]=True
    clean[couch_192]=True
    clean[table_193]=True
    clean[curtain_197]=True
    clean[curtain_198]=True
    clean[curtain_199]=True
    clean[orchid_200]=True
    clean[photoframe_210]=True
    clean[television_216]=True
    clean[light_217]=True
    clean[powersocket_218]=True
    clean[bedroom_220]=True
    clean[floor_222]=True
    clean[floor_223]=True
    clean[floor_224]=True
    clean[ceiling_226]=True
    clean[ceiling_229]=True
    clean[wall_230]=True
    clean[wall_231]=True
    clean[wall_232]=True
    clean[door_234]=True
    clean[ceilinglamp_235]=True
    clean[tablelamp_236]=True
    clean[photoframe_246]=True
    clean[light_258]=True
    clean[powersocket_259]=True
    clean[bookshelf_260]=True
    clean[desk_261]=True
    clean[nightstand_262]=True
    clean[bed_264]=True
    clean[bathroom_265]=True
    clean[wall_267]=True
    clean[wall_268]=True
    clean[wall_269]=True
    clean[wall_271]=True
    clean[floor_272]=True
    clean[floor_274]=True
    clean[floor_275]=True
    clean[ceiling_279]=True
    clean[ceiling_280]=True
    clean[ceiling_284]=True
    clean[doorjamb_285]=True
    clean[door_286]=True
    clean[ceilinglamp_288]=True
    clean[walllamp_289]=True
    clean[walllamp_290]=True
    clean[walllamp_291]=True
    clean[bathtub_297]=True
    clean[wallshelf_301]=True
    clean[toilet_302]=True
    clean[shower_303]=True
    clean[curtain_304]=True
    clean[bathroom_counter_306]=True
    clean[faucet_308]=True
    clean[light_325]=True
    clean[bedroom_327]=True
    clean[floor_330]=True
    clean[floor_334]=True
    clean[floor_336]=True
    clean[floor_337]=True
    clean[wall_340]=True
    clean[wall_341]=True
    clean[wall_342]=True
    clean[wall_343]=True
    clean[wall_344]=True
    clean[wall_345]=True
    clean[ceiling_347]=True
    clean[ceiling_348]=True
    clean[ceiling_349]=True
    clean[ceiling_351]=True
    clean[ceiling_354]=True
    clean[ceiling_355]=True
    clean[doorjamb_356]=True
    clean[ceilinglamp_357]=True
    clean[tablelamp_358]=True
    clean[tablelamp_359]=True
    clean[trashcan_360]=True
    clean[photoframe_361]=True
    clean[bookshelf_372]=True
    clean[nightstand_373]=True
    clean[desk_375]=True
    clean[bed_376]=True
    clean[dresser_377]=True
    clean[filing_cabinet_378]=True
    clean[computer_379]=True
    clean[mousepad_381]=True
    clean[cpuscreen_383]=True
    clean[light_384]=True
    clean[curtain_390]=True
    clean[curtain_391]=True
    clean[curtain_392]=True
    clean[food_orange_2008]=True
    plugged[computer_2110]=True
    plugged[light_49]=True
    plugged[fridge_140]=True
    plugged[oven_141]=True
    plugged[dishwasher_143]=True
    plugged[toaster_144]=True
    plugged[coffe_maker_147]=True
    plugged[microwave_149]=True
    plugged[television_216]=True
    plugged[light_217]=True
    plugged[light_258]=True
    plugged[light_325]=True
    plugged[computer_379]=True
    plugged[light_384]=True
    unplugged[washing_machine_2041]=True
    is_room[dining_room_1]=True
    is_room[home_office_161]=True
    is_room[bedroom_220]=True
    is_room[bathroom_265]=True
    is_room[bedroom_327]=True
    #states_end

    #char_states
    standing[char]=True
    sitting[char]=False
    lying[char]=False
    sleeping[char]=False
    has_a_free_hand[char]=True
    #char_states_end

    #char
    close_char[char,floor_15]=True
    close_char[char,kitchen_counter_128]=True
    inside_char[char,dining_room_1]=True
    #char_end

    #properties
    surfaces[chair_2118]=True
    surfaces[cutting_board_2080]=True
    surfaces[cd_player_2084]=True
    surfaces[dvd_player_2085]=True
    surfaces[stove_2090]=True
    surfaces[ironing_board_2099]=True
    surfaces[plate_2105]=True
    surfaces[floor_12]=True
    surfaces[floor_13]=True
    surfaces[floor_14]=True
    surfaces[floor_15]=True
    surfaces[floor_16]=True
    surfaces[floor_17]=True
    surfaces[floor_18]=True
    surfaces[floor_19]=True
    surfaces[floor_20]=True
    surfaces[floor_21]=True
    surfaces[floor_22]=True
    surfaces[floor_23]=True
    surfaces[floor_24]=True
    surfaces[mat_114]=True
    surfaces[mat_115]=True
    surfaces[bench_122]=True
    surfaces[table_123]=True
    surfaces[bench_124]=True
    surfaces[bench_125]=True
    surfaces[bench_126]=True
    surfaces[table_127]=True
    surfaces[kitchen_counter_128]=True
    surfaces[kitchen_counter_129]=True
    surfaces[kitchen_counter_132]=True
    surfaces[tvstand_135]=True
    surfaces[bookshelf_136]=True
    surfaces[bookshelf_137]=True
    surfaces[chair_138]=True
    surfaces[tray_142]=True
    surfaces[floor_162]=True
    surfaces[floor_163]=True
    surfaces[floor_164]=True
    surfaces[floor_165]=True
    surfaces[floor_166]=True
    surfaces[floor_167]=True
    surfaces[floor_168]=True
    surfaces[tvstand_186]=True
    surfaces[bookshelf_188]=True
    surfaces[bookshelf_189]=True
    surfaces[couch_192]=True
    surfaces[table_193]=True
    surfaces[mat_201]=True
    surfaces[floor_221]=True
    surfaces[floor_222]=True
    surfaces[floor_223]=True
    surfaces[floor_224]=True
    surfaces[floor_225]=True
    surfaces[mat_237]=True
    surfaces[bookshelf_260]=True
    surfaces[desk_261]=True
    surfaces[nightstand_262]=True
    surfaces[chair_263]=True
    surfaces[bed_264]=True
    surfaces[floor_272]=True
    surfaces[floor_273]=True
    surfaces[floor_274]=True
    surfaces[floor_275]=True
    surfaces[floor_276]=True
    surfaces[floor_277]=True
    surfaces[floor_278]=True
    surfaces[mat_292]=True
    surfaces[towel_rack_298]=True
    surfaces[towel_rack_299]=True
    surfaces[towel_rack_300]=True
    surfaces[bathroom_cabinet_305]=True
    surfaces[bathroom_counter_306]=True
    surfaces[floor_328]=True
    surfaces[floor_329]=True
    surfaces[floor_330]=True
    surfaces[floor_331]=True
    surfaces[floor_332]=True
    surfaces[floor_333]=True
    surfaces[floor_334]=True
    surfaces[floor_335]=True
    surfaces[floor_336]=True
    surfaces[floor_337]=True
    surfaces[bookshelf_372]=True
    surfaces[nightstand_373]=True
    surfaces[chair_374]=True
    surfaces[desk_375]=True
    surfaces[bed_376]=True
    surfaces[filing_cabinet_378]=True
    surfaces[mousepad_381]=True
    surfaces[mat_386]=True
    surfaces[dvd_player_2000]=True
    surfaces[stereo_2007]=True
    grabbable[keyboard_2111]=True
    grabbable[mouse_2112]=True
    grabbable[clothes_pants_2113]=True
    grabbable[clothes_shirt_2114]=True
    grabbable[clothes_socks_2115]=True
    grabbable[clothes_skirt_2116]=True
    grabbable[iron_2117]=True
    grabbable[chair_2118]=True
    grabbable[basket_for_clothes_2040]=True
    grabbable[food_steak_2042]=True
    grabbable[food_apple_2043]=True
    grabbable[food_bacon_2044]=True
    grabbable[food_banana_2045]=True
    grabbable[food_cake_2046]=True
    grabbable[food_carrot_2047]=True
    grabbable[food_cereal_2048]=True
    grabbable[food_cheese_2049]=True
    grabbable[food_chicken_2050]=True
    grabbable[food_dessert_2051]=True
    grabbable[food_donut_2052]=True
    grabbable[food_egg_2053]=True
    grabbable[food_fish_2054]=True
    grabbable[food_food_2055]=True
    grabbable[food_fruit_2056]=True
    grabbable[food_hamburger_2057]=True
    grabbable[food_ice_cream_2058]=True
    grabbable[food_jam_2059]=True
    grabbable[food_kiwi_2060]=True
    grabbable[food_lemon_2061]=True
    grabbable[food_noodles_2062]=True
    grabbable[food_oatmeal_2063]=True
    grabbable[food_peanut_butter_2064]=True
    grabbable[food_pizza_2065]=True
    grabbable[food_potato_2066]=True
    grabbable[food_rice_2067]=True
    grabbable[food_salt_2068]=True
    grabbable[food_snack_2069]=True
    grabbable[food_sugar_2070]=True
    grabbable[food_turkey_2071]=True
    grabbable[food_vegetable_2072]=True
    grabbable[dry_pasta_2073]=True
    grabbable[milk_2074]=True
    grabbable[clothes_dress_2075]=True
    grabbable[clothes_hat_2076]=True
    grabbable[clothes_gloves_2077]=True
    grabbable[clothes_jacket_2078]=True
    grabbable[clothes_scarf_2079]=True
    grabbable[cutting_board_2080]=True
    grabbable[remote_control_2081]=True
    grabbable[cat_2082]=True
    grabbable[towel_2083]=True
    grabbable[cd_player_2084]=True
    grabbable[dvd_player_2085]=True
    grabbable[headset_2086]=True
    grabbable[cup_2087]=True
    grabbable[cup_2088]=True
    grabbable[cup_2089]=True
    grabbable[book_2091]=True
    grabbable[book_2092]=True
    grabbable[pot_2093]=True
    grabbable[vacuum_cleaner_2094]=True
    grabbable[bowl_2095]=True
    grabbable[bowl_2096]=True
    grabbable[bowl_2097]=True
    grabbable[cleaning_solution_2098]=True
    grabbable[cd_2100]=True
    grabbable[sauce_2101]=True
    grabbable[oil_2102]=True
    grabbable[fork_2103]=True
    grabbable[fork_2104]=True
    grabbable[plate_2105]=True
    grabbable[spectacles_2106]=True
    grabbable[fryingpan_2107]=True
    grabbable[detergent_2108]=True
    grabbable[phone_47]=True
    grabbable[pot_54]=True
    grabbable[mat_114]=True
    grabbable[mat_115]=True
    grabbable[drawing_118]=True
    grabbable[chair_138]=True
    grabbable[tray_142]=True
    grabbable[pillow_195]=True
    grabbable[drawing_196]=True
    grabbable[mat_201]=True
    grabbable[mat_237]=True
    grabbable[drawing_238]=True
    grabbable[pillow_239]=True
    grabbable[pillow_240]=True
    grabbable[chair_263]=True
    grabbable[mat_292]=True
    grabbable[drawing_296]=True
    grabbable[towel_rack_298]=True
    grabbable[towel_rack_299]=True
    grabbable[towel_rack_300]=True
    grabbable[pillow_368]=True
    grabbable[pillow_370]=True
    grabbable[chair_374]=True
    grabbable[mouse_380]=True
    grabbable[keyboard_382]=True
    grabbable[mat_386]=True
    grabbable[drawing_387]=True
    grabbable[drawing_388]=True
    grabbable[drawing_389]=True
    grabbable[dvd_player_2000]=True
    grabbable[shoes_2001]=True
    grabbable[alcohol_2002]=True
    grabbable[mouse_2003]=True
    grabbable[coin_2004]=True
    grabbable[oil_2005]=True
    grabbable[cup_2006]=True
    grabbable[stereo_2007]=True
    grabbable[food_orange_2008]=True
    grabbable[bills_2009]=True
    grabbable[novel_2010]=True
    grabbable[homework_2011]=True
    grabbable[needle_2012]=True
    grabbable[glue_2013]=True
    grabbable[napkin_2014]=True
    grabbable[laptop_2015]=True
    grabbable[food_bread_2016]=True
    grabbable[tea_bag_2017]=True
    grabbable[food_butter_2018]=True
    grabbable[video_game_controller_2019]=True
    grabbable[crayon_2020]=True
    grabbable[dough_2021]=True
    grabbable[clothes_underwear_2022]=True
    grabbable[box_2023]=True
    grabbable[needle_2024]=True
    grabbable[laser_pointer_2025]=True
    grabbable[food_onion_2026]=True
    grabbable[console_2027]=True
    grabbable[tape_2028]=True
    grabbable[after_shave_2029]=True
    grabbable[crayon_2030]=True
    grabbable[stamp_2031]=True
    grabbable[blender_2032]=True
    grabbable[check_2033]=True
    grabbable[juice_2034]=True
    grabbable[coffee_filter_2035]=True
    grabbable[knife_2036]=True
    grabbable[soap_2037]=True
    grabbable[soap_2038]=True
    grabbable[pajamas_2039]=True
    sittable[chair_2118]=True
    sittable[mat_114]=True
    sittable[mat_115]=True
    sittable[bench_122]=True
    sittable[bench_124]=True
    sittable[bench_125]=True
    sittable[bench_126]=True
    sittable[chair_138]=True
    sittable[couch_192]=True
    sittable[mat_201]=True
    sittable[mat_237]=True
    sittable[chair_263]=True
    sittable[bed_264]=True
    sittable[mat_292]=True
    sittable[bathtub_297]=True
    sittable[toilet_302]=True
    sittable[chair_374]=True
    sittable[bed_376]=True
    sittable[mat_386]=True
    lieable[mat_114]=True
    lieable[mat_115]=True
    lieable[bench_122]=True
    lieable[bench_124]=True
    lieable[bench_125]=True
    lieable[bench_126]=True
    lieable[couch_192]=True
    lieable[mat_201]=True
    lieable[mat_237]=True
    lieable[bed_264]=True
    lieable[mat_292]=True
    lieable[bathtub_297]=True
    lieable[bed_376]=True
    lieable[mat_386]=True
    hangable[clothes_pants_2113]=True
    hangable[clothes_shirt_2114]=True
    hangable[clothes_socks_2115]=True
    hangable[clothes_skirt_2116]=True
    hangable[clothes_dress_2075]=True
    hangable[clothes_hat_2076]=True
    hangable[clothes_gloves_2077]=True
    hangable[clothes_jacket_2078]=True
    hangable[clothes_scarf_2079]=True
    hangable[clothes_underwear_2022]=True
    drinkable[milk_2074]=True
    drinkable[oil_2102]=True
    drinkable[alcohol_2002]=True
    drinkable[oil_2005]=True
    drinkable[juice_2034]=True
    eatable[food_steak_2042]=True
    eatable[food_apple_2043]=True
    eatable[food_bacon_2044]=True
    eatable[food_banana_2045]=True
    eatable[food_cake_2046]=True
    eatable[food_carrot_2047]=True
    eatable[food_cereal_2048]=True
    eatable[food_cheese_2049]=True
    eatable[food_chicken_2050]=True
    eatable[food_dessert_2051]=True
    eatable[food_egg_2053]=True
    eatable[food_fish_2054]=True
    eatable[food_food_2055]=True
    eatable[food_fruit_2056]=True
    eatable[food_hamburger_2057]=True
    eatable[food_jam_2059]=True
    eatable[food_kiwi_2060]=True
    eatable[food_lemon_2061]=True
    eatable[food_noodles_2062]=True
    eatable[food_oatmeal_2063]=True
    eatable[food_peanut_butter_2064]=True
    eatable[food_pizza_2065]=True
    eatable[food_potato_2066]=True
    eatable[food_rice_2067]=True
    eatable[food_salt_2068]=True
    eatable[food_snack_2069]=True
    eatable[food_sugar_2070]=True
    eatable[food_turkey_2071]=True
    eatable[food_vegetable_2072]=True
    eatable[food_orange_2008]=True
    eatable[food_bread_2016]=True
    eatable[food_onion_2026]=True
    recipient[washing_machine_2041]=True
    recipient[cup_2087]=True
    recipient[cup_2088]=True
    recipient[cup_2089]=True
    recipient[pot_2093]=True
    recipient[bowl_2095]=True
    recipient[bowl_2096]=True
    recipient[bowl_2097]=True
    recipient[plate_2105]=True
    recipient[fryingpan_2107]=True
    recipient[pot_54]=True
    recipient[sink_133]=True
    recipient[coffe_maker_147]=True
    recipient[sink_307]=True
    recipient[cup_2006]=True
    recipient[box_2023]=True
    recipient[blender_2032]=True
    cuttable[food_steak_2042]=True
    cuttable[food_apple_2043]=True
    cuttable[food_bacon_2044]=True
    cuttable[food_banana_2045]=True
    cuttable[food_cake_2046]=True
    cuttable[food_carrot_2047]=True
    cuttable[food_cheese_2049]=True
    cuttable[food_chicken_2050]=True
    cuttable[food_dessert_2051]=True
    cuttable[food_egg_2053]=True
    cuttable[food_fish_2054]=True
    cuttable[food_food_2055]=True
    cuttable[food_fruit_2056]=True
    cuttable[food_hamburger_2057]=True
    cuttable[food_kiwi_2060]=True
    cuttable[food_lemon_2061]=True
    cuttable[food_pizza_2065]=True
    cuttable[food_potato_2066]=True
    cuttable[food_turkey_2071]=True
    cuttable[food_vegetable_2072]=True
    cuttable[book_2091]=True
    cuttable[book_2092]=True
    cuttable[drawing_118]=True
    cuttable[drawing_196]=True
    cuttable[drawing_238]=True
    cuttable[drawing_296]=True
    cuttable[drawing_387]=True
    cuttable[drawing_388]=True
    cuttable[drawing_389]=True
    cuttable[food_orange_2008]=True
    cuttable[bills_2009]=True
    cuttable[novel_2010]=True
    cuttable[food_bread_2016]=True
    cuttable[food_onion_2026]=True
    pourable[food_cereal_2048]=True
    pourable[food_rice_2067]=True
    pourable[food_salt_2068]=True
    pourable[food_sugar_2070]=True
    pourable[milk_2074]=True
    pourable[cup_2087]=True
    pourable[cup_2088]=True
    pourable[cup_2089]=True
    pourable[cleaning_solution_2098]=True
    pourable[sauce_2101]=True
    pourable[oil_2102]=True
    pourable[detergent_2108]=True
    pourable[alcohol_2002]=True
    pourable[oil_2005]=True
    pourable[cup_2006]=True
    pourable[after_shave_2029]=True
    pourable[blender_2032]=True
    pourable[juice_2034]=True
    can_open[basket_for_clothes_2040]=True
    can_open[washing_machine_2041]=True
    can_open[food_cereal_2048]=True
    can_open[food_jam_2059]=True
    can_open[milk_2074]=True
    can_open[cd_player_2084]=True
    can_open[dvd_player_2085]=True
    can_open[stove_2090]=True
    can_open[book_2091]=True
    can_open[book_2092]=True
    can_open[pot_2093]=True
    can_open[window_2109]=True
    can_open[door_38]=True
    can_open[window_40]=True
    can_open[pot_54]=True
    can_open[curtain_119]=True
    can_open[curtain_120]=True
    can_open[curtain_121]=True
    can_open[cupboard_130]=True
    can_open[cupboard_131]=True
    can_open[bookshelf_136]=True
    can_open[bookshelf_137]=True
    can_open[fridge_140]=True
    can_open[oven_141]=True
    can_open[dishwasher_143]=True
    can_open[coffe_maker_147]=True
    can_open[microwave_149]=True
    can_open[window_181]=True
    can_open[bookshelf_188]=True
    can_open[bookshelf_189]=True
    can_open[curtain_197]=True
    can_open[curtain_198]=True
    can_open[curtain_199]=True
    can_open[door_234]=True
    can_open[bookshelf_260]=True
    can_open[nightstand_262]=True
    can_open[door_286]=True
    can_open[window_287]=True
    can_open[curtain_293]=True
    can_open[curtain_294]=True
    can_open[toilet_302]=True
    can_open[curtain_304]=True
    can_open[bathroom_cabinet_305]=True
    can_open[window_346]=True
    can_open[trashcan_360]=True
    can_open[bookshelf_372]=True
    can_open[nightstand_373]=True
    can_open[dresser_377]=True
    can_open[filing_cabinet_378]=True
    can_open[curtain_390]=True
    can_open[curtain_391]=True
    can_open[curtain_392]=True
    can_open[dvd_player_2000]=True
    can_open[stereo_2007]=True
    can_open[novel_2010]=True
    can_open[box_2023]=True
    can_open[console_2027]=True
    can_open[after_shave_2029]=True
    can_open[blender_2032]=True
    has_switch[iron_2117]=True
    has_switch[washing_machine_2041]=True
    has_switch[remote_control_2081]=True
    has_switch[cd_player_2084]=True
    has_switch[dvd_player_2085]=True
    has_switch[stove_2090]=True
    has_switch[vacuum_cleaner_2094]=True
    has_switch[computer_2110]=True
    has_switch[phone_47]=True
    has_switch[light_49]=True
    has_switch[faucet_134]=True
    has_switch[fridge_140]=True
    has_switch[oven_141]=True
    has_switch[dishwasher_143]=True
    has_switch[toaster_144]=True
    has_switch[coffe_maker_147]=True
    has_switch[microwave_149]=True
    has_switch[television_216]=True
    has_switch[light_217]=True
    has_switch[tablelamp_236]=True
    has_switch[light_258]=True
    has_switch[faucet_308]=True
    has_switch[light_325]=True
    has_switch[tablelamp_358]=True
    has_switch[tablelamp_359]=True
    has_switch[computer_379]=True
    has_switch[light_384]=True
    has_switch[dvd_player_2000]=True
    has_switch[stereo_2007]=True
    has_switch[laptop_2015]=True
    has_switch[video_game_controller_2019]=True
    has_switch[laser_pointer_2025]=True
    has_switch[console_2027]=True
    has_switch[blender_2032]=True
    containers[basket_for_clothes_2040]=True
    containers[washing_machine_2041]=True
    containers[cd_player_2084]=True
    containers[stove_2090]=True
    containers[pot_2093]=True
    containers[fryingpan_2107]=True
    containers[pot_54]=True
    containers[cupboard_130]=True
    containers[cupboard_131]=True
    containers[sink_133]=True
    containers[bookshelf_136]=True
    containers[bookshelf_137]=True
    containers[fridge_140]=True
    containers[oven_141]=True
    containers[dishwasher_143]=True
    containers[toaster_144]=True
    containers[coffe_maker_147]=True
    containers[microwave_149]=True
    containers[bookshelf_188]=True
    containers[bookshelf_189]=True
    containers[bookshelf_260]=True
    containers[nightstand_262]=True
    containers[toilet_302]=True
    containers[bathroom_cabinet_305]=True
    containers[sink_307]=True
    containers[trashcan_360]=True
    containers[bookshelf_372]=True
    containers[nightstand_373]=True
    containers[dresser_377]=True
    containers[filing_cabinet_378]=True
    containers[box_2023]=True
    has_plug[keyboard_2111]=True
    has_plug[mouse_2112]=True
    has_plug[iron_2117]=True
    has_plug[washing_machine_2041]=True
    has_plug[cd_player_2084]=True
    has_plug[dvd_player_2085]=True
    has_plug[vacuum_cleaner_2094]=True
    has_plug[phone_47]=True
    has_plug[light_49]=True
    has_plug[fridge_140]=True
    has_plug[oven_141]=True
    has_plug[toaster_144]=True
    has_plug[coffe_maker_147]=True
    has_plug[microwave_149]=True
    has_plug[television_216]=True
    has_plug[light_217]=True
    has_plug[light_258]=True
    has_plug[light_325]=True
    has_plug[mouse_380]=True
    has_plug[keyboard_382]=True
    has_plug[light_384]=True
    has_plug[dvd_player_2000]=True
    has_plug[mouse_2003]=True
    has_plug[stereo_2007]=True
    has_plug[laptop_2015]=True
    has_plug[video_game_controller_2019]=True
    has_plug[console_2027]=True
    has_plug[blender_2032]=True
    readable[book_2091]=True
    readable[book_2092]=True
    readable[bills_2009]=True
    readable[novel_2010]=True
    readable[homework_2011]=True
    readable[check_2033]=True
    lookable[computer_2110]=True
    lookable[drawing_118]=True
    lookable[drawing_196]=True
    lookable[television_216]=True
    lookable[drawing_238]=True
    lookable[drawing_296]=True
    lookable[computer_379]=True
    lookable[drawing_387]=True
    lookable[drawing_388]=True
    lookable[drawing_389]=True
    lookable[laptop_2015]=True
    is_clothes[clothes_pants_2113]=True
    is_clothes[clothes_shirt_2114]=True
    is_clothes[clothes_socks_2115]=True
    is_clothes[clothes_skirt_2116]=True
    is_clothes[clothes_dress_2075]=True
    is_clothes[clothes_hat_2076]=True
    is_clothes[clothes_gloves_2077]=True
    is_clothes[clothes_jacket_2078]=True
    is_clothes[clothes_scarf_2079]=True
    is_clothes[headset_2086]=True
    is_clothes[spectacles_2106]=True
    is_clothes[shoes_2001]=True
    is_clothes[clothes_underwear_2022]=True
    is_clothes[pajamas_2039]=True
    is_food[food_steak_2042]=True
    is_food[food_apple_2043]=True
    is_food[food_bacon_2044]=True
    is_food[food_banana_2045]=True
    is_food[food_cake_2046]=True
    is_food[food_carrot_2047]=True
    is_food[food_cereal_2048]=True
    is_food[food_cheese_2049]=True
    is_food[food_chicken_2050]=True
    is_food[food_dessert_2051]=True
    is_food[food_donut_2052]=True
    is_food[food_egg_2053]=True
    is_food[food_fish_2054]=True
    is_food[food_food_2055]=True
    is_food[food_fruit_2056]=True
    is_food[food_hamburger_2057]=True
    is_food[food_ice_cream_2058]=True
    is_food[food_jam_2059]=True
    is_food[food_kiwi_2060]=True
    is_food[food_lemon_2061]=True
    is_food[food_noodles_2062]=True
    is_food[food_oatmeal_2063]=True
    is_food[food_peanut_butter_2064]=True
    is_food[food_pizza_2065]=True
    is_food[food_potato_2066]=True
    is_food[food_rice_2067]=True
    is_food[food_salt_2068]=True
    is_food[food_snack_2069]=True
    is_food[food_sugar_2070]=True
    is_food[food_turkey_2071]=True
    is_food[food_vegetable_2072]=True
    is_food[food_orange_2008]=True
    is_food[food_bread_2016]=True
    is_food[food_butter_2018]=True
    is_food[food_onion_2026]=True
    cover_object[towel_2083]=True
    cover_object[curtain_119]=True
    cover_object[curtain_120]=True
    cover_object[curtain_121]=True
    cover_object[curtain_197]=True
    cover_object[curtain_198]=True
    cover_object[curtain_199]=True
    cover_object[curtain_293]=True
    cover_object[curtain_294]=True
    cover_object[curtain_304]=True
    cover_object[curtain_390]=True
    cover_object[curtain_391]=True
    cover_object[curtain_392]=True
    cover_object[napkin_2014]=True
    cover_object[box_2023]=True
    has_paper[book_2091]=True
    has_paper[book_2092]=True
    has_paper[drawing_118]=True
    has_paper[drawing_196]=True
    has_paper[drawing_238]=True
    has_paper[drawing_296]=True
    has_paper[drawing_387]=True
    has_paper[drawing_388]=True
    has_paper[drawing_389]=True
    has_paper[bills_2009]=True
    has_paper[novel_2010]=True
    has_paper[homework_2011]=True
    has_paper[napkin_2014]=True
    has_paper[check_2033]=True
    has_paper[coffee_filter_2035]=True
    movable[keyboard_2111]=True
    movable[mouse_2112]=True
    movable[clothes_pants_2113]=True
    movable[clothes_shirt_2114]=True
    movable[clothes_socks_2115]=True
    movable[clothes_skirt_2116]=True
    movable[iron_2117]=True
    movable[chair_2118]=True
    movable[basket_for_clothes_2040]=True
    movable[food_steak_2042]=True
    movable[food_apple_2043]=True
    movable[food_bacon_2044]=True
    movable[food_banana_2045]=True
    movable[food_cake_2046]=True
    movable[food_carrot_2047]=True
    movable[food_cereal_2048]=True
    movable[food_cheese_2049]=True
    movable[food_chicken_2050]=True
    movable[food_dessert_2051]=True
    movable[food_donut_2052]=True
    movable[food_egg_2053]=True
    movable[food_fish_2054]=True
    movable[food_food_2055]=True
    movable[food_fruit_2056]=True
    movable[food_hamburger_2057]=True
    movable[food_ice_cream_2058]=True
    movable[food_jam_2059]=True
    movable[food_kiwi_2060]=True
    movable[food_lemon_2061]=True
    movable[food_noodles_2062]=True
    movable[food_oatmeal_2063]=True
    movable[food_peanut_butter_2064]=True
    movable[food_pizza_2065]=True
    movable[food_potato_2066]=True
    movable[food_rice_2067]=True
    movable[food_salt_2068]=True
    movable[food_snack_2069]=True
    movable[food_sugar_2070]=True
    movable[food_turkey_2071]=True
    movable[food_vegetable_2072]=True
    movable[dry_pasta_2073]=True
    movable[milk_2074]=True
    movable[clothes_dress_2075]=True
    movable[clothes_hat_2076]=True
    movable[clothes_gloves_2077]=True
    movable[clothes_jacket_2078]=True
    movable[clothes_scarf_2079]=True
    movable[cutting_board_2080]=True
    movable[remote_control_2081]=True
    movable[cat_2082]=True
    movable[towel_2083]=True
    movable[cd_player_2084]=True
    movable[dvd_player_2085]=True
    movable[headset_2086]=True
    movable[cup_2087]=True
    movable[cup_2088]=True
    movable[cup_2089]=True
    movable[book_2091]=True
    movable[book_2092]=True
    movable[pot_2093]=True
    movable[vacuum_cleaner_2094]=True
    movable[bowl_2095]=True
    movable[bowl_2096]=True
    movable[bowl_2097]=True
    movable[cleaning_solution_2098]=True
    movable[ironing_board_2099]=True
    movable[cd_2100]=True
    movable[sauce_2101]=True
    movable[oil_2102]=True
    movable[fork_2103]=True
    movable[fork_2104]=True
    movable[plate_2105]=True
    movable[spectacles_2106]=True
    movable[fryingpan_2107]=True
    movable[detergent_2108]=True
    movable[phone_47]=True
    movable[pot_54]=True
    movable[mat_114]=True
    movable[mat_115]=True
    movable[drawing_118]=True
    movable[curtain_119]=True
    movable[curtain_120]=True
    movable[curtain_121]=True
    movable[bench_122]=True
    movable[table_123]=True
    movable[bench_124]=True
    movable[bench_125]=True
    movable[bench_126]=True
    movable[table_127]=True
    movable[chair_138]=True
    movable[tray_142]=True
    movable[toaster_144]=True
    movable[coffe_maker_147]=True
    movable[couch_192]=True
    movable[table_193]=True
    movable[pillow_195]=True
    movable[drawing_196]=True
    movable[curtain_197]=True
    movable[curtain_198]=True
    movable[curtain_199]=True
    movable[mat_201]=True
    movable[mat_237]=True
    movable[drawing_238]=True
    movable[pillow_239]=True
    movable[pillow_240]=True
    movable[desk_261]=True
    movable[chair_263]=True
    movable[mat_292]=True
    movable[curtain_293]=True
    movable[curtain_294]=True
    movable[drawing_296]=True
    movable[towel_rack_298]=True
    movable[towel_rack_299]=True
    movable[towel_rack_300]=True
    movable[curtain_304]=True
    movable[trashcan_360]=True
    movable[pillow_368]=True
    movable[pillow_370]=True
    movable[chair_374]=True
    movable[desk_375]=True
    movable[mouse_380]=True
    movable[mousepad_381]=True
    movable[keyboard_382]=True
    movable[mat_386]=True
    movable[drawing_387]=True
    movable[drawing_388]=True
    movable[drawing_389]=True
    movable[curtain_390]=True
    movable[curtain_391]=True
    movable[curtain_392]=True
    movable[dvd_player_2000]=True
    movable[shoes_2001]=True
    movable[alcohol_2002]=True
    movable[mouse_2003]=True
    movable[coin_2004]=True
    movable[oil_2005]=True
    movable[cup_2006]=True
    movable[stereo_2007]=True
    movable[food_orange_2008]=True
    movable[bills_2009]=True
    movable[novel_2010]=True
    movable[homework_2011]=True
    movable[needle_2012]=True
    movable[glue_2013]=True
    movable[napkin_2014]=True
    movable[laptop_2015]=True
    movable[food_bread_2016]=True
    movable[tea_bag_2017]=True
    movable[food_butter_2018]=True
    movable[video_game_controller_2019]=True
    movable[crayon_2020]=True
    movable[dough_2021]=True
    movable[clothes_underwear_2022]=True
    movable[box_2023]=True
    movable[needle_2024]=True
    movable[laser_pointer_2025]=True
    movable[food_onion_2026]=True
    movable[console_2027]=True
    movable[tape_2028]=True
    movable[after_shave_2029]=True
    movable[crayon_2030]=True
    movable[stamp_2031]=True
    movable[blender_2032]=True
    movable[check_2033]=True
    movable[juice_2034]=True
    movable[coffee_filter_2035]=True
    movable[knife_2036]=True
    movable[soap_2037]=True
    movable[soap_2038]=True
    movable[pajamas_2039]=True
    cream[food_cheese_2049]=True
    cream[food_ice_cream_2058]=True
    cream[food_jam_2059]=True
    cream[food_peanut_butter_2064]=True
    cream[sauce_2101]=True
    cream[glue_2013]=True
    cream[food_butter_2018]=True
    cream[dough_2021]=True
    cream[after_shave_2029]=True
    cream[soap_2037]=True
    cream[soap_2038]=True
    #properties_end

    #relations
    on[cutting_board_2080,kitchen_counter_128]=True
    on[stove_2090,kitchen_counter_129]=True
    on[spectacles_2106,kitchen_counter_128]=True
    on[computer_2110,table_193]=True
    on[ceiling_25,wall_5]=True
    on[ceiling_27,wall_6]=True
    on[ceiling_34,wall_7]=True
    on[ceiling_36,wall_11]=True
    on[door_38,floor_336]=True
    on[knifeblock_52,wall_2]=True
    on[orchid_117,tvstand_135]=True
    on[table_123,floor_17]=True
    on[table_127,floor_20]=True
    on[kitchen_counter_128,floor_15]=True
    on[faucet_134,kitchen_counter_132]=True
    on[tvstand_135,floor_19]=True
    on[bookshelf_136,floor_12]=True
    on[bookshelf_136,floor_13]=True
    on[bookshelf_137,floor_24]=True
    on[fridge_140,floor_22]=True
    on[dishwasher_143,floor_21]=True
    on[toaster_144,kitchen_counter_129]=True
    on[coffe_maker_147,kitchen_counter_129]=True
    on[microwave_149,kitchen_counter_132]=True
    on[wall_170,floor_164]=True
    on[ceiling_175,wall_169]=True
    on[ceiling_176,wall_171]=True
    on[ceiling_179,wall_170]=True
    on[ceiling_180,wall_174]=True
    on[tvstand_186,floor_162]=True
    on[tvstand_186,floor_163]=True
    on[bookshelf_188,floor_165]=True
    on[bookshelf_189,floor_167]=True
    on[orchid_200,table_193]=True
    on[photoframe_210,wallshelf_187]=True
    on[television_216,tvstand_186]=True
    on[ceiling_226,wall_233]=True
    on[ceiling_227,wall_231]=True
    on[ceiling_228,wall_232]=True
    on[ceiling_229,wall_230]=True
    on[door_234,floor_165]=True
    on[door_234,floor_224]=True
    on[tablelamp_236,nightstand_262]=True
    on[bookshelf_260,floor_221]=True
    on[bookshelf_260,floor_222]=True
    on[desk_261,floor_223]=True
    on[nightstand_262,floor_221]=True
    on[nightstand_262,floor_222]=True
    on[ceiling_279,wall_269]=True
    on[ceiling_281,wall_268]=True
    on[ceiling_282,wall_267]=True
    on[ceiling_284,wall_266]=True
    on[doorjamb_285,floor_337]=True
    on[door_286,floor_337]=True
    on[bathroom_cabinet_305,wall_269]=True
    on[faucet_308,bathroom_counter_306]=True
    on[ceiling_347,wall_341]=True
    on[ceiling_349,wall_342]=True
    on[ceiling_353,wall_343]=True
    on[ceiling_355,wall_345]=True
    on[tablelamp_358,bed_376]=True
    on[tablelamp_359,nightstand_373]=True
    on[trashcan_360,floor_328]=True
    on[trashcan_360,floor_329]=True
    on[photoframe_361,bookshelf_372]=True
    on[bookshelf_372,floor_331]=True
    on[nightstand_373,floor_330]=True
    on[desk_375,floor_337]=True
    on[bed_376,floor_330]=True
    on[filing_cabinet_378,floor_335]=True
    on[mousepad_381,desk_375]=True
    on[cpuscreen_383,desk_375]=True
    on[food_orange_2008,kitchen_counter_128]=True
    inside[washing_machine_2041,bathroom_265]=True
    inside[stove_2090,dining_room_1]=True
    inside[ironing_board_2099,bedroom_220]=True
    inside[window_2109,dining_room_1]=True
    inside[computer_2110,home_office_161]=True
    inside[wall_2,dining_room_1]=True
    inside[wall_3,dining_room_1]=True
    inside[wall_4,dining_room_1]=True
    inside[wall_5,dining_room_1]=True
    inside[wall_6,dining_room_1]=True
    inside[wall_7,dining_room_1]=True
    inside[wall_8,dining_room_1]=True
    inside[wall_9,dining_room_1]=True
    inside[wall_10,dining_room_1]=True
    inside[wall_11,dining_room_1]=True
    inside[floor_12,dining_room_1]=True
    inside[floor_13,dining_room_1]=True
    inside[floor_14,dining_room_1]=True
    inside[floor_15,dining_room_1]=True
    inside[floor_16,dining_room_1]=True
    inside[floor_17,dining_room_1]=True
    inside[floor_18,dining_room_1]=True
    inside[floor_19,dining_room_1]=True
    inside[floor_20,dining_room_1]=True
    inside[floor_21,dining_room_1]=True
    inside[floor_22,dining_room_1]=True
    inside[floor_23,dining_room_1]=True
    inside[floor_24,dining_room_1]=True
    inside[ceiling_25,dining_room_1]=True
    inside[ceiling_26,dining_room_1]=True
    inside[ceiling_27,dining_room_1]=True
    inside[ceiling_28,dining_room_1]=True
    inside[ceiling_29,dining_room_1]=True
    inside[ceiling_30,dining_room_1]=True
    inside[ceiling_31,dining_room_1]=True
    inside[ceiling_32,dining_room_1]=True
    inside[ceiling_33,dining_room_1]=True
    inside[ceiling_34,dining_room_1]=True
    inside[ceiling_35,dining_room_1]=True
    inside[ceiling_36,dining_room_1]=True
    inside[doorjamb_37,dining_room_1]=True
    inside[door_38,dining_room_1]=True
    inside[doorjamb_39,dining_room_1]=True
    inside[window_40,dining_room_1]=True
    inside[ceilinglamp_41,dining_room_1]=True
    inside[ceilinglamp_42,dining_room_1]=True
    inside[ceilinglamp_43,dining_room_1]=True
    inside[walllamp_44,dining_room_1]=True
    inside[walllamp_45,dining_room_1]=True
    inside[walllamp_46,dining_room_1]=True
    inside[powersocket_48,dining_room_1]=True
    inside[light_49,dining_room_1]=True
    inside[knifeblock_52,dining_room_1]=True
    inside[photoframe_102,dining_room_1]=True
    inside[photoframe_102,bookshelf_137]=True
    inside[orchid_117,dining_room_1]=True
    inside[curtain_119,dining_room_1]=True
    inside[curtain_119,curtain_120]=True
    inside[curtain_120,dining_room_1]=True
    inside[curtain_120,curtain_119]=True
    inside[curtain_121,dining_room_1]=True
    inside[bench_122,dining_room_1]=True
    inside[table_123,dining_room_1]=True
    inside[bench_124,dining_room_1]=True
    inside[bench_125,dining_room_1]=True
    inside[bench_126,dining_room_1]=True
    inside[table_127,dining_room_1]=True
    inside[kitchen_counter_128,dining_room_1]=True
    inside[kitchen_counter_129,dining_room_1]=True
    inside[cupboard_130,dining_room_1]=True
    inside[cupboard_131,dining_room_1]=True
    inside[kitchen_counter_132,dining_room_1]=True
    inside[sink_133,dining_room_1]=True
    inside[sink_133,kitchen_counter_132]=True
    inside[faucet_134,dining_room_1]=True
    inside[tvstand_135,dining_room_1]=True
    inside[bookshelf_136,dining_room_1]=True
    inside[bookshelf_137,dining_room_1]=True
    inside[stovefan_139,dining_room_1]=True
    inside[fridge_140,dining_room_1]=True
    inside[oven_141,dining_room_1]=True
    inside[dishwasher_143,dining_room_1]=True
    inside[toaster_144,dining_room_1]=True
    inside[coffe_maker_147,dining_room_1]=True
    inside[microwave_149,dining_room_1]=True
    inside[floor_162,home_office_161]=True
    inside[floor_163,home_office_161]=True
    inside[floor_164,home_office_161]=True
    inside[floor_165,home_office_161]=True
    inside[floor_166,home_office_161]=True
    inside[floor_167,home_office_161]=True
    inside[floor_168,home_office_161]=True
    inside[wall_169,home_office_161]=True
    inside[wall_170,home_office_161]=True
    inside[wall_171,home_office_161]=True
    inside[wall_172,home_office_161]=True
    inside[wall_173,home_office_161]=True
    inside[wall_174,home_office_161]=True
    inside[ceiling_175,home_office_161]=True
    inside[ceiling_176,home_office_161]=True
    inside[ceiling_177,home_office_161]=True
    inside[ceiling_178,home_office_161]=True
    inside[ceiling_179,home_office_161]=True
    inside[ceiling_180,home_office_161]=True
    inside[window_181,home_office_161]=True
    inside[doorjamb_182,home_office_161]=True
    inside[walllamp_183,home_office_161]=True
    inside[walllamp_184,home_office_161]=True
    inside[ceilinglamp_185,home_office_161]=True
    inside[tvstand_186,home_office_161]=True
    inside[wallshelf_187,home_office_161]=True
    inside[bookshelf_188,home_office_161]=True
    inside[bookshelf_189,home_office_161]=True
    inside[wallshelf_190,home_office_161]=True
    inside[wallshelf_191,home_office_161]=True
    inside[couch_192,home_office_161]=True
    inside[table_193,home_office_161]=True
    inside[curtain_197,home_office_161]=True
    inside[curtain_197,curtain_198]=True
    inside[curtain_198,home_office_161]=True
    inside[curtain_198,curtain_197]=True
    inside[curtain_199,home_office_161]=True
    inside[orchid_200,home_office_161]=True
    inside[photoframe_210,home_office_161]=True
    inside[television_216,home_office_161]=True
    inside[light_217,home_office_161]=True
    inside[powersocket_218,home_office_161]=True
    inside[floor_221,bedroom_220]=True
    inside[floor_222,bedroom_220]=True
    inside[floor_223,bedroom_220]=True
    inside[floor_224,bedroom_220]=True
    inside[floor_225,bedroom_220]=True
    inside[ceiling_226,bedroom_220]=True
    inside[ceiling_227,bedroom_220]=True
    inside[ceiling_228,bedroom_220]=True
    inside[ceiling_229,bedroom_220]=True
    inside[wall_230,bedroom_220]=True
    inside[wall_231,bedroom_220]=True
    inside[wall_232,bedroom_220]=True
    inside[wall_233,bedroom_220]=True
    inside[door_234,bedroom_220]=True
    inside[ceilinglamp_235,bedroom_220]=True
    inside[tablelamp_236,bedroom_220]=True
    inside[photoframe_246,bedroom_220]=True
    inside[photoframe_246,bookshelf_260]=True
    inside[light_258,bedroom_220]=True
    inside[powersocket_259,bedroom_220]=True
    inside[bookshelf_260,bedroom_220]=True
    inside[desk_261,bedroom_220]=True
    inside[nightstand_262,bedroom_220]=True
    inside[bed_264,bedroom_220]=True
    inside[wall_266,bathroom_265]=True
    inside[wall_267,bathroom_265]=True
    inside[wall_268,bathroom_265]=True
    inside[wall_269,bathroom_265]=True
    inside[wall_270,bathroom_265]=True
    inside[wall_271,bathroom_265]=True
    inside[floor_272,bathroom_265]=True
    inside[floor_273,bathroom_265]=True
    inside[floor_274,bathroom_265]=True
    inside[floor_275,bathroom_265]=True
    inside[floor_276,bathroom_265]=True
    inside[floor_277,bathroom_265]=True
    inside[floor_278,bathroom_265]=True
    inside[ceiling_279,bathroom_265]=True
    inside[ceiling_280,bathroom_265]=True
    inside[ceiling_281,bathroom_265]=True
    inside[ceiling_282,bathroom_265]=True
    inside[ceiling_283,bathroom_265]=True
    inside[ceiling_284,bathroom_265]=True
    inside[doorjamb_285,bathroom_265]=True
    inside[door_286,bathroom_265]=True
    inside[window_287,bathroom_265]=True
    inside[ceilinglamp_288,bathroom_265]=True
    inside[walllamp_289,bathroom_265]=True
    inside[walllamp_290,bathroom_265]=True
    inside[walllamp_291,bathroom_265]=True
    inside[curtain_293,bathroom_265]=True
    inside[curtain_293,curtain_294]=True
    inside[curtain_294,bathroom_265]=True
    inside[curtain_294,curtain_293]=True
    inside[bathtub_297,bathroom_265]=True
    inside[wallshelf_301,bathroom_265]=True
    inside[toilet_302,bathroom_265]=True
    inside[shower_303,bathroom_265]=True
    inside[curtain_304,bathroom_265]=True
    inside[curtain_304,shower_303]=True
    inside[bathroom_cabinet_305,bathroom_265]=True
    inside[bathroom_counter_306,bathroom_265]=True
    inside[sink_307,bathroom_265]=True
    inside[sink_307,bathroom_counter_306]=True
    inside[faucet_308,bathroom_265]=True
    inside[light_325,bathroom_265]=True
    inside[floor_328,bedroom_327]=True
    inside[floor_329,bedroom_327]=True
    inside[floor_330,bedroom_327]=True
    inside[floor_331,bedroom_327]=True
    inside[floor_332,bedroom_327]=True
    inside[floor_333,bedroom_327]=True
    inside[floor_334,bedroom_327]=True
    inside[floor_335,bedroom_327]=True
    inside[floor_336,bedroom_327]=True
    inside[floor_337,bedroom_327]=True
    inside[wall_338,bedroom_327]=True
    inside[wall_339,bedroom_327]=True
    inside[wall_340,bedroom_327]=True
    inside[wall_341,bedroom_327]=True
    inside[wall_342,bedroom_327]=True
    inside[wall_343,bedroom_327]=True
    inside[wall_344,bedroom_327]=True
    inside[wall_345,bedroom_327]=True
    inside[window_346,bedroom_327]=True
    inside[ceiling_347,bedroom_327]=True
    inside[ceiling_348,bedroom_327]=True
    inside[ceiling_349,bedroom_327]=True
    inside[ceiling_350,bedroom_327]=True
    inside[ceiling_351,bedroom_327]=True
    inside[ceiling_352,bedroom_327]=True
    inside[ceiling_353,bedroom_327]=True
    inside[ceiling_354,bedroom_327]=True
    inside[ceiling_355,bedroom_327]=True
    inside[doorjamb_356,bedroom_327]=True
    inside[ceilinglamp_357,bedroom_327]=True
    inside[tablelamp_358,bedroom_327]=True
    inside[tablelamp_359,bedroom_327]=True
    inside[trashcan_360,bedroom_327]=True
    inside[photoframe_361,bedroom_327]=True
    inside[bookshelf_372,bedroom_327]=True
    inside[nightstand_373,bedroom_327]=True
    inside[desk_375,bedroom_327]=True
    inside[bed_376,bedroom_327]=True
    inside[dresser_377,bedroom_327]=True
    inside[filing_cabinet_378,bedroom_327]=True
    inside[computer_379,bedroom_327]=True
    inside[mousepad_381,bedroom_327]=True
    inside[cpuscreen_383,bedroom_327]=True
    inside[light_384,bedroom_327]=True
    inside[curtain_390,bedroom_327]=True
    inside[curtain_390,curtain_391]=True
    inside[curtain_391,bedroom_327]=True
    inside[curtain_391,curtain_390]=True
    inside[curtain_392,bedroom_327]=True
    between[doorjamb_37,dining_room_1]=True
    between[doorjamb_37,home_office_161]=True
    between[door_38,dining_room_1]=True
    between[door_38,bedroom_327]=True
    between[door_234,home_office_161]=True
    between[door_234,bedroom_220]=True
    between[door_286,bathroom_265]=True
    between[door_286,bedroom_327]=True
    close[washing_machine_2041,window_287]=True
    close[washing_machine_2041,bathtub_297]=True
    close[cutting_board_2080,kitchen_counter_128]=True
    close[stove_2090,kitchen_counter_129]=True
    close[ironing_board_2099,bedroom_220]=True
    close[spectacles_2106,kitchen_counter_128]=True
    close[window_2109,dining_room_1]=True
    close[computer_2110,table_193]=True
    close[dining_room_1,window_2109]=True
    close[wall_2,wall_6]=True
    close[wall_2,wall_8]=True
    close[wall_2,floor_16]=True
    close[wall_2,ceiling_28]=True
    close[wall_2,walllamp_45]=True
    close[wall_2,walllamp_46]=True
    close[wall_2,knifeblock_52]=True
    close[wall_2,kitchen_counter_129]=True
    close[wall_2,cupboard_130]=True
    close[wall_2,cupboard_131]=True
    close[wall_2,kitchen_counter_132]=True
    close[wall_2,sink_133]=True
    close[wall_2,faucet_134]=True
    close[wall_2,stovefan_139]=True
    close[wall_2,oven_141]=True
    close[wall_2,microwave_149]=True
    close[wall_3,wall_5]=True
    close[wall_3,wall_6]=True
    close[wall_3,floor_14]=True
    close[wall_3,ceiling_26]=True
    close[wall_3,doorjamb_37]=True
    close[wall_3,powersocket_48]=True
    close[wall_3,light_49]=True
    close[wall_3,floor_166]=True
    close[wall_3,wall_171]=True
    close[wall_3,wall_172]=True
    close[wall_3,ceiling_176]=True
    close[wall_3,walllamp_183]=True
    close[wall_3,bookshelf_189]=True
    close[wall_3,light_217]=True
    close[wall_3,powersocket_218]=True
    close[wall_3,wall_268]=True
    close[wall_3,toilet_302]=True
    close[wall_4,wall_7]=True
    close[wall_4,wall_11]=True
    close[wall_4,floor_23]=True
    close[wall_4,ceiling_35]=True
    close[wall_4,doorjamb_39]=True
    close[wall_4,window_40]=True
    close[wall_4,ceilinglamp_43]=True
    close[wall_4,curtain_119]=True
    close[wall_4,curtain_120]=True
    close[wall_4,curtain_121]=True
    close[wall_5,wall_3]=True
    close[wall_5,wall_10]=True
    close[wall_5,floor_12]=True
    close[wall_5,floor_13]=True
    close[wall_5,floor_14]=True
    close[wall_5,floor_18]=True
    close[wall_5,ceiling_25]=True
    close[wall_5,ceiling_26]=True
    close[wall_5,ceiling_30]=True
    close[wall_5,doorjamb_37]=True
    close[wall_5,door_38]=True
    close[wall_5,ceilinglamp_41]=True
    close[wall_5,powersocket_48]=True
    close[wall_5,light_49]=True
    close[wall_5,table_123]=True
    close[wall_5,bench_124]=True
    close[wall_5,bookshelf_136]=True
    close[wall_5,walllamp_183]=True
    close[wall_5,wall_268]=True
    close[wall_5,wall_271]=True
    close[wall_5,floor_277]=True
    close[wall_5,ceiling_281]=True
    close[wall_5,doorjamb_285]=True
    close[wall_5,door_286]=True
    close[wall_5,toilet_302]=True
    close[wall_5,floor_337]=True
    close[wall_5,wall_344]=True
    close[wall_5,wall_345]=True
    close[wall_5,ceiling_355]=True
    close[wall_5,doorjamb_356]=True
    close[wall_5,desk_375]=True
    close[wall_5,computer_379]=True
    close[wall_5,mousepad_381]=True
    close[wall_5,cpuscreen_383]=True
    close[wall_6,wall_2]=True
    close[wall_6,wall_3]=True
    close[wall_6,floor_14]=True
    close[wall_6,floor_15]=True
    close[wall_6,floor_16]=True
    close[wall_6,ceiling_26]=True
    close[wall_6,ceiling_27]=True
    close[wall_6,ceiling_28]=True
    close[wall_6,doorjamb_37]=True
    close[wall_6,ceilinglamp_41]=True
    close[wall_6,walllamp_45]=True
    close[wall_6,knifeblock_52]=True
    close[wall_6,bench_122]=True
    close[wall_6,kitchen_counter_128]=True
    close[wall_6,cupboard_130]=True
    close[wall_6,kitchen_counter_132]=True
    close[wall_6,sink_133]=True
    close[wall_6,faucet_134]=True
    close[wall_6,microwave_149]=True
    close[wall_6,floor_167]=True
    close[wall_6,wall_172]=True
    close[wall_6,ceiling_177]=True
    close[wall_6,bookshelf_188]=True
    close[wall_6,bookshelf_189]=True
    close[wall_6,light_217]=True
    close[wall_6,powersocket_218]=True
    close[wall_7,wall_4]=True
    close[wall_7,wall_8]=True
    close[wall_7,floor_21]=True
    close[wall_7,floor_22]=True
    close[wall_7,floor_23]=True
    close[wall_7,ceiling_33]=True
    close[wall_7,ceiling_34]=True
    close[wall_7,ceiling_35]=True
    close[wall_7,window_40]=True
    close[wall_7,ceilinglamp_43]=True
    close[wall_7,walllamp_44]=True
    close[wall_7,curtain_119]=True
    close[wall_7,curtain_120]=True
    close[wall_7,bench_126]=True
    close[wall_7,kitchen_counter_129]=True
    close[wall_7,cupboard_131]=True
    close[wall_7,fridge_140]=True
    close[wall_7,dishwasher_143]=True
    close[wall_7,toaster_144]=True
    close[wall_7,coffe_maker_147]=True
    close[wall_8,wall_2]=True
    close[wall_8,wall_7]=True
    close[wall_8,floor_21]=True
    close[wall_8,ceiling_33]=True
    close[wall_8,walllamp_44]=True
    close[wall_8,walllamp_46]=True
    close[wall_8,knifeblock_52]=True
    close[wall_8,kitchen_counter_129]=True
    close[wall_8,cupboard_131]=True
    close[wall_8,stovefan_139]=True
    close[wall_8,fridge_140]=True
    close[wall_8,oven_141]=True
    close[wall_8,dishwasher_143]=True
    close[wall_8,toaster_144]=True
    close[wall_8,coffe_maker_147]=True
    close[wall_9,wall_10]=True
    close[wall_9,wall_11]=True
    close[wall_9,floor_19]=True
    close[wall_9,ceiling_31]=True
    close[wall_9,door_38]=True
    close[wall_9,orchid_117]=True
    close[wall_9,tvstand_135]=True
    close[wall_9,bookshelf_137]=True
    close[wall_9,floor_335]=True
    close[wall_9,wall_343]=True
    close[wall_9,wall_344]=True
    close[wall_9,ceiling_353]=True
    close[wall_9,doorjamb_356]=True
    close[wall_9,filing_cabinet_378]=True
    close[wall_9,light_384]=True
    close[wall_10,wall_5]=True
    close[wall_10,wall_9]=True
    close[wall_10,floor_18]=True
    close[wall_10,ceiling_30]=True
    close[wall_10,door_38]=True
    close[wall_10,orchid_117]=True
    close[wall_10,tvstand_135]=True
    close[wall_10,bookshelf_136]=True
    close[wall_10,floor_336]=True
    close[wall_10,wall_343]=True
    close[wall_10,wall_344]=True
    close[wall_10,wall_345]=True
    close[wall_10,ceiling_354]=True
    close[wall_10,doorjamb_356]=True
    close[wall_10,desk_375]=True
    close[wall_10,computer_379]=True
    close[wall_10,mousepad_381]=True
    close[wall_10,cpuscreen_383]=True
    close[wall_10,light_384]=True
    close[wall_11,wall_4]=True
    close[wall_11,wall_9]=True
    close[wall_11,floor_19]=True
    close[wall_11,floor_23]=True
    close[wall_11,floor_24]=True
    close[wall_11,ceiling_31]=True
    close[wall_11,ceiling_35]=True
    close[wall_11,ceiling_36]=True
    close[wall_11,doorjamb_39]=True
    close[wall_11,window_40]=True
    close[wall_11,ceilinglamp_43]=True
    close[wall_11,photoframe_102]=True
    close[wall_11,curtain_121]=True
    close[wall_11,bench_125]=True
    close[wall_11,table_127]=True
    close[wall_11,bookshelf_137]=True
    close[wall_11,filing_cabinet_378]=True
    close[floor_12,wall_5]=True
    close[floor_12,floor_13]=True
    close[floor_12,floor_14]=True
    close[floor_12,floor_18]=True
    close[floor_12,door_38]=True
    close[floor_12,powersocket_48]=True
    close[floor_12,light_49]=True
    close[floor_12,table_123]=True
    close[floor_12,bench_124]=True
    close[floor_12,bookshelf_136]=True
    close[floor_12,wall_268]=True
    close[floor_12,floor_277]=True
    close[floor_12,door_286]=True
    close[floor_12,toilet_302]=True
    close[floor_12,floor_337]=True
    close[floor_12,wall_345]=True
    close[floor_12,desk_375]=True
    close[floor_12,computer_379]=True
    close[floor_12,mousepad_381]=True
    close[floor_12,cpuscreen_383]=True
    close[floor_13,wall_5]=True
    close[floor_13,floor_12]=True
    close[floor_13,floor_14]=True
    close[floor_13,floor_18]=True
    close[floor_13,door_38]=True
    close[floor_13,powersocket_48]=True
    close[floor_13,light_49]=True
    close[floor_13,table_123]=True
    close[floor_13,bench_124]=True
    close[floor_13,bookshelf_136]=True
    close[floor_13,wall_268]=True
    close[floor_13,floor_277]=True
    close[floor_13,door_286]=True
    close[floor_13,toilet_302]=True
    close[floor_13,floor_337]=True
    close[floor_13,wall_345]=True
    close[floor_13,desk_375]=True
    close[floor_13,computer_379]=True
    close[floor_13,mousepad_381]=True
    close[floor_13,cpuscreen_383]=True
    close[floor_14,wall_3]=True
    close[floor_14,wall_5]=True
    close[floor_14,wall_6]=True
    close[floor_14,floor_12]=True
    close[floor_14,floor_13]=True
    close[floor_14,floor_15]=True
    close[floor_14,floor_17]=True
    close[floor_14,doorjamb_37]=True
    close[floor_14,powersocket_48]=True
    close[floor_14,light_49]=True
    close[floor_14,bench_122]=True
    close[floor_14,table_123]=True
    close[floor_14,bench_124]=True
    close[floor_14,floor_166]=True
    close[floor_14,wall_171]=True
    close[floor_14,bookshelf_189]=True
    close[floor_14,light_217]=True
    close[floor_14,powersocket_218]=True
    close[floor_14,toilet_302]=True
    close[floor_15,wall_6]=True
    close[floor_15,floor_14]=True
    close[floor_15,floor_16]=True
    close[floor_15,bench_122]=True
    close[floor_15,kitchen_counter_128]=True
    close[floor_15,kitchen_counter_132]=True
    close[floor_15,sink_133]=True
    close[floor_15,faucet_134]=True
    close[floor_15,microwave_149]=True
    close[floor_15,floor_167]=True
    close[floor_15,wall_172]=True
    close[floor_15,bookshelf_188]=True
    close[floor_15,bookshelf_189]=True
    close[floor_15,light_217]=True
    close[floor_15,powersocket_218]=True
    close[floor_16,wall_2]=True
    close[floor_16,wall_6]=True
    close[floor_16,floor_15]=True
    close[floor_16,floor_17]=True
    close[floor_16,floor_21]=True
    close[floor_16,knifeblock_52]=True
    close[floor_16,bench_122]=True
    close[floor_16,kitchen_counter_129]=True
    close[floor_16,kitchen_counter_132]=True
    close[floor_16,sink_133]=True
    close[floor_16,faucet_134]=True
    close[floor_16,oven_141]=True
    close[floor_17,floor_14]=True
    close[floor_17,floor_16]=True
    close[floor_17,floor_18]=True
    close[floor_17,floor_20]=True
    close[floor_17,bench_122]=True
    close[floor_17,table_123]=True
    close[floor_17,bench_124]=True
    close[floor_18,wall_5]=True
    close[floor_18,wall_10]=True
    close[floor_18,floor_12]=True
    close[floor_18,floor_13]=True
    close[floor_18,floor_17]=True
    close[floor_18,floor_19]=True
    close[floor_18,door_38]=True
    close[floor_18,orchid_117]=True
    close[floor_18,table_123]=True
    close[floor_18,bench_124]=True
    close[floor_18,tvstand_135]=True
    close[floor_18,bookshelf_136]=True
    close[floor_18,floor_336]=True
    close[floor_18,wall_344]=True
    close[floor_18,doorjamb_356]=True
    close[floor_18,desk_375]=True
    close[floor_18,computer_379]=True
    close[floor_18,mousepad_381]=True
    close[floor_18,cpuscreen_383]=True
    close[floor_18,light_384]=True
    close[floor_19,wall_9]=True
    close[floor_19,wall_11]=True
    close[floor_19,floor_18]=True
    close[floor_19,floor_20]=True
    close[floor_19,floor_24]=True
    close[floor_19,door_38]=True
    close[floor_19,orchid_117]=True
    close[floor_19,bench_125]=True
    close[floor_19,table_127]=True
    close[floor_19,tvstand_135]=True
    close[floor_19,bookshelf_137]=True
    close[floor_19,floor_335]=True
    close[floor_19,wall_343]=True
    close[floor_19,light_384]=True
    close[floor_20,floor_17]=True
    close[floor_20,floor_19]=True
    close[floor_20,floor_21]=True
    close[floor_20,floor_23]=True
    close[floor_20,bench_125]=True
    close[floor_20,bench_126]=True
    close[floor_20,table_127]=True
    close[floor_21,wall_7]=True
    close[floor_21,wall_8]=True
    close[floor_21,floor_16]=True
    close[floor_21,floor_20]=True
    close[floor_21,floor_22]=True
    close[floor_21,bench_126]=True
    close[floor_21,kitchen_counter_129]=True
    close[floor_21,oven_141]=True
    close[floor_21,dishwasher_143]=True
    close[floor_21,toaster_144]=True
    close[floor_21,coffe_maker_147]=True
    close[floor_22,wall_7]=True
    close[floor_22,floor_21]=True
    close[floor_22,floor_23]=True
    close[floor_22,bench_126]=True
    close[floor_22,kitchen_counter_129]=True
    close[floor_22,fridge_140]=True
    close[floor_22,dishwasher_143]=True
    close[floor_22,toaster_144]=True
    close[floor_23,wall_4]=True
    close[floor_23,wall_7]=True
    close[floor_23,wall_11]=True
    close[floor_23,floor_20]=True
    close[floor_23,floor_22]=True
    close[floor_23,floor_24]=True
    close[floor_23,window_40]=True
    close[floor_23,curtain_119]=True
    close[floor_23,curtain_120]=True
    close[floor_23,curtain_121]=True
    close[floor_23,bench_125]=True
    close[floor_23,bench_126]=True
    close[floor_23,table_127]=True
    close[floor_24,wall_11]=True
    close[floor_24,floor_19]=True
    close[floor_24,floor_23]=True
    close[floor_24,doorjamb_39]=True
    close[floor_24,photoframe_102]=True
    close[floor_24,bench_125]=True
    close[floor_24,table_127]=True
    close[floor_24,bookshelf_137]=True
    close[ceiling_25,wall_5]=True
    close[ceiling_25,ceiling_26]=True
    close[ceiling_25,ceiling_30]=True
    close[ceiling_25,ceilinglamp_41]=True
    close[ceiling_25,light_49]=True
    close[ceiling_25,bookshelf_136]=True
    close[ceiling_25,walllamp_183]=True
    close[ceiling_25,wall_268]=True
    close[ceiling_25,ceiling_281]=True
    close[ceiling_25,wall_345]=True
    close[ceiling_25,ceiling_355]=True
    close[ceiling_25,cpuscreen_383]=True
    close[ceiling_26,wall_3]=True
    close[ceiling_26,wall_5]=True
    close[ceiling_26,wall_6]=True
    close[ceiling_26,ceiling_25]=True
    close[ceiling_26,ceiling_27]=True
    close[ceiling_26,ceiling_29]=True
    close[ceiling_26,doorjamb_37]=True
    close[ceiling_26,ceilinglamp_41]=True
    close[ceiling_26,light_49]=True
    close[ceiling_26,wall_171]=True
    close[ceiling_26,ceiling_176]=True
    close[ceiling_26,walllamp_183]=True
    close[ceiling_26,light_217]=True
    close[ceiling_27,wall_6]=True
    close[ceiling_27,ceiling_26]=True
    close[ceiling_27,ceiling_28]=True
    close[ceiling_27,ceilinglamp_41]=True
    close[ceiling_27,walllamp_45]=True
    close[ceiling_27,knifeblock_52]=True
    close[ceiling_27,kitchen_counter_128]=True
    close[ceiling_27,cupboard_130]=True
    close[ceiling_27,faucet_134]=True
    close[ceiling_27,microwave_149]=True
    close[ceiling_27,wall_172]=True
    close[ceiling_27,ceiling_177]=True
    close[ceiling_27,bookshelf_189]=True
    close[ceiling_27,light_217]=True
    close[ceiling_28,wall_2]=True
    close[ceiling_28,wall_6]=True
    close[ceiling_28,ceiling_27]=True
    close[ceiling_28,ceiling_29]=True
    close[ceiling_28,ceiling_33]=True
    close[ceiling_28,ceilinglamp_41]=True
    close[ceiling_28,ceilinglamp_42]=True
    close[ceiling_28,walllamp_45]=True
    close[ceiling_28,walllamp_46]=True
    close[ceiling_28,knifeblock_52]=True
    close[ceiling_28,cupboard_130]=True
    close[ceiling_28,faucet_134]=True
    close[ceiling_28,stovefan_139]=True
    close[ceiling_29,ceiling_26]=True
    close[ceiling_29,ceiling_28]=True
    close[ceiling_29,ceiling_30]=True
    close[ceiling_29,ceiling_32]=True
    close[ceiling_29,ceilinglamp_41]=True
    close[ceiling_29,ceilinglamp_42]=True
    close[ceiling_30,wall_5]=True
    close[ceiling_30,wall_10]=True
    close[ceiling_30,ceiling_25]=True
    close[ceiling_30,ceiling_29]=True
    close[ceiling_30,ceiling_31]=True
    close[ceiling_30,ceilinglamp_41]=True
    close[ceiling_30,ceilinglamp_42]=True
    close[ceiling_30,bookshelf_136]=True
    close[ceiling_30,wall_344]=True
    close[ceiling_30,ceiling_354]=True
    close[ceiling_30,doorjamb_356]=True
    close[ceiling_30,cpuscreen_383]=True
    close[ceiling_30,light_384]=True
    close[ceiling_31,wall_9]=True
    close[ceiling_31,wall_11]=True
    close[ceiling_31,ceiling_30]=True
    close[ceiling_31,ceiling_32]=True
    close[ceiling_31,ceiling_36]=True
    close[ceiling_31,ceilinglamp_42]=True
    close[ceiling_31,bookshelf_137]=True
    close[ceiling_31,wall_343]=True
    close[ceiling_31,ceiling_353]=True
    close[ceiling_31,light_384]=True
    close[ceiling_32,ceiling_29]=True
    close[ceiling_32,ceiling_31]=True
    close[ceiling_32,ceiling_33]=True
    close[ceiling_32,ceiling_35]=True
    close[ceiling_32,ceilinglamp_42]=True
    close[ceiling_32,ceilinglamp_43]=True
    close[ceiling_33,wall_7]=True
    close[ceiling_33,wall_8]=True
    close[ceiling_33,ceiling_28]=True
    close[ceiling_33,ceiling_32]=True
    close[ceiling_33,ceiling_34]=True
    close[ceiling_33,ceilinglamp_42]=True
    close[ceiling_33,walllamp_44]=True
    close[ceiling_33,walllamp_46]=True
    close[ceiling_33,cupboard_131]=True
    close[ceiling_33,stovefan_139]=True
    close[ceiling_33,toaster_144]=True
    close[ceiling_33,coffe_maker_147]=True
    close[ceiling_34,wall_7]=True
    close[ceiling_34,ceiling_33]=True
    close[ceiling_34,ceiling_35]=True
    close[ceiling_34,ceilinglamp_43]=True
    close[ceiling_34,walllamp_44]=True
    close[ceiling_34,curtain_119]=True
    close[ceiling_34,curtain_120]=True
    close[ceiling_34,cupboard_131]=True
    close[ceiling_34,fridge_140]=True
    close[ceiling_34,toaster_144]=True
    close[ceiling_34,coffe_maker_147]=True
    close[ceiling_35,wall_4]=True
    close[ceiling_35,wall_7]=True
    close[ceiling_35,wall_11]=True
    close[ceiling_35,ceiling_32]=True
    close[ceiling_35,ceiling_34]=True
    close[ceiling_35,ceiling_36]=True
    close[ceiling_35,window_40]=True
    close[ceiling_35,ceilinglamp_43]=True
    close[ceiling_35,curtain_119]=True
    close[ceiling_35,curtain_120]=True
    close[ceiling_35,curtain_121]=True
    close[ceiling_36,wall_11]=True
    close[ceiling_36,ceiling_31]=True
    close[ceiling_36,ceiling_35]=True
    close[ceiling_36,doorjamb_39]=True
    close[ceiling_36,ceilinglamp_43]=True
    close[ceiling_36,photoframe_102]=True
    close[ceiling_36,curtain_121]=True
    close[ceiling_36,bookshelf_137]=True
    close[doorjamb_37,wall_3]=True
    close[doorjamb_37,wall_5]=True
    close[doorjamb_37,wall_6]=True
    close[doorjamb_37,floor_14]=True
    close[doorjamb_37,ceiling_26]=True
    close[doorjamb_37,powersocket_48]=True
    close[doorjamb_37,light_49]=True
    close[doorjamb_37,floor_166]=True
    close[doorjamb_37,wall_171]=True
    close[doorjamb_37,wall_172]=True
    close[doorjamb_37,ceiling_176]=True
    close[doorjamb_37,walllamp_183]=True
    close[doorjamb_37,bookshelf_189]=True
    close[doorjamb_37,light_217]=True
    close[doorjamb_37,powersocket_218]=True
    close[doorjamb_37,wall_268]=True
    close[door_38,wall_5]=True
    close[door_38,wall_9]=True
    close[door_38,wall_10]=True
    close[door_38,floor_12]=True
    close[door_38,floor_13]=True
    close[door_38,floor_18]=True
    close[door_38,floor_19]=True
    close[door_38,orchid_117]=True
    close[door_38,bookshelf_136]=True
    close[door_38,floor_335]=True
    close[door_38,floor_336]=True
    close[door_38,floor_337]=True
    close[door_38,wall_343]=True
    close[door_38,wall_344]=True
    close[door_38,wall_345]=True
    close[door_38,doorjamb_356]=True
    close[door_38,desk_375]=True
    close[door_38,mousepad_381]=True
    close[door_38,cpuscreen_383]=True
    close[door_38,light_384]=True
    close[doorjamb_39,wall_4]=True
    close[doorjamb_39,wall_11]=True
    close[doorjamb_39,floor_24]=True
    close[doorjamb_39,ceiling_36]=True
    close[doorjamb_39,window_40]=True
    close[doorjamb_39,photoframe_102]=True
    close[doorjamb_39,curtain_121]=True
    close[doorjamb_39,bookshelf_137]=True
    close[window_40,wall_4]=True
    close[window_40,wall_7]=True
    close[window_40,wall_11]=True
    close[window_40,floor_23]=True
    close[window_40,ceiling_35]=True
    close[window_40,doorjamb_39]=True
    close[window_40,ceilinglamp_43]=True
    close[window_40,curtain_119]=True
    close[window_40,curtain_120]=True
    close[window_40,curtain_121]=True
    close[ceilinglamp_41,wall_5]=True
    close[ceilinglamp_41,wall_6]=True
    close[ceilinglamp_41,ceiling_25]=True
    close[ceilinglamp_41,ceiling_26]=True
    close[ceilinglamp_41,ceiling_27]=True
    close[ceilinglamp_41,ceiling_28]=True
    close[ceilinglamp_41,ceiling_29]=True
    close[ceilinglamp_41,ceiling_30]=True
    close[ceilinglamp_41,table_123]=True
    close[ceilinglamp_42,ceiling_28]=True
    close[ceilinglamp_42,ceiling_29]=True
    close[ceilinglamp_42,ceiling_30]=True
    close[ceilinglamp_42,ceiling_31]=True
    close[ceilinglamp_42,ceiling_32]=True
    close[ceilinglamp_42,ceiling_33]=True
    close[ceilinglamp_43,wall_4]=True
    close[ceilinglamp_43,wall_7]=True
    close[ceilinglamp_43,wall_11]=True
    close[ceilinglamp_43,ceiling_32]=True
    close[ceilinglamp_43,ceiling_34]=True
    close[ceilinglamp_43,ceiling_35]=True
    close[ceilinglamp_43,ceiling_36]=True
    close[ceilinglamp_43,window_40]=True
    close[ceilinglamp_43,curtain_119]=True
    close[ceilinglamp_43,curtain_120]=True
    close[ceilinglamp_43,curtain_121]=True
    close[walllamp_44,wall_7]=True
    close[walllamp_44,wall_8]=True
    close[walllamp_44,ceiling_33]=True
    close[walllamp_44,ceiling_34]=True
    close[walllamp_44,kitchen_counter_129]=True
    close[walllamp_44,cupboard_131]=True
    close[walllamp_44,dishwasher_143]=True
    close[walllamp_44,toaster_144]=True
    close[walllamp_44,coffe_maker_147]=True
    close[walllamp_45,wall_2]=True
    close[walllamp_45,wall_6]=True
    close[walllamp_45,ceiling_27]=True
    close[walllamp_45,ceiling_28]=True
    close[walllamp_45,knifeblock_52]=True
    close[walllamp_45,cupboard_130]=True
    close[walllamp_45,kitchen_counter_132]=True
    close[walllamp_45,sink_133]=True
    close[walllamp_45,faucet_134]=True
    close[walllamp_45,microwave_149]=True
    close[walllamp_46,wall_2]=True
    close[walllamp_46,wall_8]=True
    close[walllamp_46,ceiling_28]=True
    close[walllamp_46,ceiling_33]=True
    close[walllamp_46,knifeblock_52]=True
    close[walllamp_46,kitchen_counter_129]=True
    close[walllamp_46,cupboard_130]=True
    close[walllamp_46,cupboard_131]=True
    close[walllamp_46,kitchen_counter_132]=True
    close[walllamp_46,stovefan_139]=True
    close[walllamp_46,oven_141]=True
    close[powersocket_48,wall_3]=True
    close[powersocket_48,wall_5]=True
    close[powersocket_48,floor_12]=True
    close[powersocket_48,floor_13]=True
    close[powersocket_48,floor_14]=True
    close[powersocket_48,doorjamb_37]=True
    close[powersocket_48,light_49]=True
    close[powersocket_48,floor_166]=True
    close[powersocket_48,wall_171]=True
    close[powersocket_48,tvstand_186]=True
    close[powersocket_48,light_217]=True
    close[powersocket_48,powersocket_218]=True
    close[powersocket_48,wall_268]=True
    close[powersocket_48,floor_277]=True
    close[powersocket_48,toilet_302]=True
    close[light_49,wall_3]=True
    close[light_49,wall_5]=True
    close[light_49,floor_12]=True
    close[light_49,floor_13]=True
    close[light_49,floor_14]=True
    close[light_49,ceiling_25]=True
    close[light_49,ceiling_26]=True
    close[light_49,doorjamb_37]=True
    close[light_49,powersocket_48]=True
    close[light_49,floor_166]=True
    close[light_49,wall_171]=True
    close[light_49,ceiling_176]=True
    close[light_49,walllamp_183]=True
    close[light_49,light_217]=True
    close[light_49,powersocket_218]=True
    close[light_49,wall_268]=True
    close[light_49,floor_277]=True
    close[light_49,toilet_302]=True
    close[knifeblock_52,wall_2]=True
    close[knifeblock_52,wall_6]=True
    close[knifeblock_52,wall_8]=True
    close[knifeblock_52,floor_16]=True
    close[knifeblock_52,ceiling_27]=True
    close[knifeblock_52,ceiling_28]=True
    close[knifeblock_52,walllamp_45]=True
    close[knifeblock_52,walllamp_46]=True
    close[knifeblock_52,cupboard_130]=True
    close[knifeblock_52,kitchen_counter_132]=True
    close[knifeblock_52,sink_133]=True
    close[knifeblock_52,faucet_134]=True
    close[knifeblock_52,stovefan_139]=True
    close[knifeblock_52,oven_141]=True
    close[photoframe_102,wall_11]=True
    close[photoframe_102,floor_24]=True
    close[photoframe_102,ceiling_36]=True
    close[photoframe_102,doorjamb_39]=True
    close[photoframe_102,bookshelf_137]=True
    close[orchid_117,wall_9]=True
    close[orchid_117,wall_10]=True
    close[orchid_117,floor_18]=True
    close[orchid_117,floor_19]=True
    close[orchid_117,door_38]=True
    close[orchid_117,tvstand_135]=True
    close[orchid_117,floor_335]=True
    close[orchid_117,floor_336]=True
    close[orchid_117,wall_343]=True
    close[orchid_117,wall_344]=True
    close[orchid_117,light_384]=True
    close[curtain_119,wall_4]=True
    close[curtain_119,wall_7]=True
    close[curtain_119,floor_23]=True
    close[curtain_119,ceiling_34]=True
    close[curtain_119,ceiling_35]=True
    close[curtain_119,window_40]=True
    close[curtain_119,ceilinglamp_43]=True
    close[curtain_119,curtain_120]=True
    close[curtain_119,curtain_121]=True
    close[curtain_120,wall_4]=True
    close[curtain_120,wall_7]=True
    close[curtain_120,floor_23]=True
    close[curtain_120,ceiling_34]=True
    close[curtain_120,ceiling_35]=True
    close[curtain_120,window_40]=True
    close[curtain_120,ceilinglamp_43]=True
    close[curtain_120,curtain_119]=True
    close[curtain_120,curtain_121]=True
    close[curtain_121,wall_4]=True
    close[curtain_121,wall_11]=True
    close[curtain_121,floor_23]=True
    close[curtain_121,ceiling_35]=True
    close[curtain_121,ceiling_36]=True
    close[curtain_121,doorjamb_39]=True
    close[curtain_121,window_40]=True
    close[curtain_121,ceilinglamp_43]=True
    close[curtain_121,curtain_119]=True
    close[curtain_121,curtain_120]=True
    close[bench_122,wall_6]=True
    close[bench_122,floor_14]=True
    close[bench_122,floor_15]=True
    close[bench_122,floor_16]=True
    close[bench_122,floor_17]=True
    close[bench_122,table_123]=True
    close[bench_122,bench_124]=True
    close[table_123,wall_5]=True
    close[table_123,floor_12]=True
    close[table_123,floor_13]=True
    close[table_123,floor_14]=True
    close[table_123,floor_17]=True
    close[table_123,floor_18]=True
    close[table_123,ceilinglamp_41]=True
    close[table_123,bench_122]=True
    close[table_123,bench_124]=True
    close[bench_124,wall_5]=True
    close[bench_124,floor_12]=True
    close[bench_124,floor_13]=True
    close[bench_124,floor_14]=True
    close[bench_124,floor_17]=True
    close[bench_124,floor_18]=True
    close[bench_124,bench_122]=True
    close[bench_124,table_123]=True
    close[bench_125,wall_11]=True
    close[bench_125,floor_19]=True
    close[bench_125,floor_20]=True
    close[bench_125,floor_23]=True
    close[bench_125,floor_24]=True
    close[bench_125,bench_126]=True
    close[bench_125,table_127]=True
    close[bench_126,wall_7]=True
    close[bench_126,floor_20]=True
    close[bench_126,floor_21]=True
    close[bench_126,floor_22]=True
    close[bench_126,floor_23]=True
    close[bench_126,bench_125]=True
    close[bench_126,table_127]=True
    close[table_127,wall_11]=True
    close[table_127,floor_19]=True
    close[table_127,floor_20]=True
    close[table_127,floor_23]=True
    close[table_127,floor_24]=True
    close[table_127,bench_125]=True
    close[table_127,bench_126]=True
    close[kitchen_counter_128,cutting_board_2080]=True
    close[kitchen_counter_128,spectacles_2106]=True
    close[kitchen_counter_128,wall_6]=True
    close[kitchen_counter_128,floor_15]=True
    close[kitchen_counter_128,ceiling_27]=True
    close[kitchen_counter_128,cupboard_130]=True
    close[kitchen_counter_128,kitchen_counter_132]=True
    close[kitchen_counter_128,sink_133]=True
    close[kitchen_counter_128,microwave_149]=True
    close[kitchen_counter_128,floor_165]=True
    close[kitchen_counter_128,floor_167]=True
    close[kitchen_counter_128,wall_172]=True
    close[kitchen_counter_128,wall_174]=True
    close[kitchen_counter_128,bookshelf_188]=True
    close[kitchen_counter_128,bookshelf_189]=True
    close[kitchen_counter_128,food_orange_2008]=True
    close[kitchen_counter_129,stove_2090]=True
    close[kitchen_counter_129,wall_2]=True
    close[kitchen_counter_129,wall_7]=True
    close[kitchen_counter_129,wall_8]=True
    close[kitchen_counter_129,floor_16]=True
    close[kitchen_counter_129,floor_21]=True
    close[kitchen_counter_129,floor_22]=True
    close[kitchen_counter_129,walllamp_44]=True
    close[kitchen_counter_129,walllamp_46]=True
    close[kitchen_counter_129,cupboard_131]=True
    close[kitchen_counter_129,stovefan_139]=True
    close[kitchen_counter_129,fridge_140]=True
    close[kitchen_counter_129,oven_141]=True
    close[kitchen_counter_129,dishwasher_143]=True
    close[kitchen_counter_129,toaster_144]=True
    close[kitchen_counter_129,coffe_maker_147]=True
    close[cupboard_130,wall_2]=True
    close[cupboard_130,wall_6]=True
    close[cupboard_130,ceiling_27]=True
    close[cupboard_130,ceiling_28]=True
    close[cupboard_130,walllamp_45]=True
    close[cupboard_130,walllamp_46]=True
    close[cupboard_130,knifeblock_52]=True
    close[cupboard_130,kitchen_counter_128]=True
    close[cupboard_130,kitchen_counter_132]=True
    close[cupboard_130,sink_133]=True
    close[cupboard_130,faucet_134]=True
    close[cupboard_130,stovefan_139]=True
    close[cupboard_130,oven_141]=True
    close[cupboard_130,microwave_149]=True
    close[cupboard_130,wall_172]=True
    close[cupboard_131,wall_2]=True
    close[cupboard_131,wall_7]=True
    close[cupboard_131,wall_8]=True
    close[cupboard_131,ceiling_33]=True
    close[cupboard_131,ceiling_34]=True
    close[cupboard_131,walllamp_44]=True
    close[cupboard_131,walllamp_46]=True
    close[cupboard_131,kitchen_counter_129]=True
    close[cupboard_131,stovefan_139]=True
    close[cupboard_131,fridge_140]=True
    close[cupboard_131,oven_141]=True
    close[cupboard_131,dishwasher_143]=True
    close[cupboard_131,toaster_144]=True
    close[cupboard_131,coffe_maker_147]=True
    close[kitchen_counter_132,wall_2]=True
    close[kitchen_counter_132,wall_6]=True
    close[kitchen_counter_132,floor_15]=True
    close[kitchen_counter_132,floor_16]=True
    close[kitchen_counter_132,walllamp_45]=True
    close[kitchen_counter_132,walllamp_46]=True
    close[kitchen_counter_132,knifeblock_52]=True
    close[kitchen_counter_132,kitchen_counter_128]=True
    close[kitchen_counter_132,cupboard_130]=True
    close[kitchen_counter_132,sink_133]=True
    close[kitchen_counter_132,faucet_134]=True
    close[kitchen_counter_132,stovefan_139]=True
    close[kitchen_counter_132,oven_141]=True
    close[kitchen_counter_132,microwave_149]=True
    close[kitchen_counter_132,wall_172]=True
    close[sink_133,wall_2]=True
    close[sink_133,wall_6]=True
    close[sink_133,floor_15]=True
    close[sink_133,floor_16]=True
    close[sink_133,walllamp_45]=True
    close[sink_133,knifeblock_52]=True
    close[sink_133,kitchen_counter_128]=True
    close[sink_133,cupboard_130]=True
    close[sink_133,kitchen_counter_132]=True
    close[sink_133,faucet_134]=True
    close[sink_133,microwave_149]=True
    close[faucet_134,wall_2]=True
    close[faucet_134,wall_6]=True
    close[faucet_134,floor_15]=True
    close[faucet_134,floor_16]=True
    close[faucet_134,ceiling_27]=True
    close[faucet_134,ceiling_28]=True
    close[faucet_134,walllamp_45]=True
    close[faucet_134,knifeblock_52]=True
    close[faucet_134,cupboard_130]=True
    close[faucet_134,kitchen_counter_132]=True
    close[faucet_134,sink_133]=True
    close[faucet_134,oven_141]=True
    close[faucet_134,microwave_149]=True
    close[tvstand_135,wall_9]=True
    close[tvstand_135,wall_10]=True
    close[tvstand_135,floor_18]=True
    close[tvstand_135,floor_19]=True
    close[tvstand_135,orchid_117]=True
    close[tvstand_135,bookshelf_137]=True
    close[tvstand_135,floor_335]=True
    close[tvstand_135,floor_336]=True
    close[tvstand_135,wall_343]=True
    close[tvstand_135,wall_344]=True
    close[tvstand_135,light_384]=True
    close[bookshelf_136,wall_5]=True
    close[bookshelf_136,wall_10]=True
    close[bookshelf_136,floor_12]=True
    close[bookshelf_136,floor_13]=True
    close[bookshelf_136,floor_18]=True
    close[bookshelf_136,ceiling_25]=True
    close[bookshelf_136,ceiling_30]=True
    close[bookshelf_136,door_38]=True
    close[bookshelf_136,doorjamb_285]=True
    close[bookshelf_136,door_286]=True
    close[bookshelf_136,floor_336]=True
    close[bookshelf_136,floor_337]=True
    close[bookshelf_136,wall_344]=True
    close[bookshelf_136,wall_345]=True
    close[bookshelf_136,ceiling_355]=True
    close[bookshelf_136,doorjamb_356]=True
    close[bookshelf_136,desk_375]=True
    close[bookshelf_136,computer_379]=True
    close[bookshelf_136,mousepad_381]=True
    close[bookshelf_136,cpuscreen_383]=True
    close[bookshelf_137,wall_9]=True
    close[bookshelf_137,wall_11]=True
    close[bookshelf_137,floor_19]=True
    close[bookshelf_137,floor_24]=True
    close[bookshelf_137,ceiling_31]=True
    close[bookshelf_137,ceiling_36]=True
    close[bookshelf_137,doorjamb_39]=True
    close[bookshelf_137,photoframe_102]=True
    close[bookshelf_137,tvstand_135]=True
    close[bookshelf_137,floor_335]=True
    close[bookshelf_137,wall_343]=True
    close[bookshelf_137,filing_cabinet_378]=True
    close[stovefan_139,wall_2]=True
    close[stovefan_139,wall_8]=True
    close[stovefan_139,ceiling_28]=True
    close[stovefan_139,ceiling_33]=True
    close[stovefan_139,walllamp_46]=True
    close[stovefan_139,knifeblock_52]=True
    close[stovefan_139,kitchen_counter_129]=True
    close[stovefan_139,cupboard_130]=True
    close[stovefan_139,cupboard_131]=True
    close[stovefan_139,kitchen_counter_132]=True
    close[stovefan_139,oven_141]=True
    close[fridge_140,wall_7]=True
    close[fridge_140,wall_8]=True
    close[fridge_140,floor_22]=True
    close[fridge_140,ceiling_34]=True
    close[fridge_140,kitchen_counter_129]=True
    close[fridge_140,cupboard_131]=True
    close[fridge_140,toaster_144]=True
    close[oven_141,wall_2]=True
    close[oven_141,wall_8]=True
    close[oven_141,floor_16]=True
    close[oven_141,floor_21]=True
    close[oven_141,walllamp_46]=True
    close[oven_141,knifeblock_52]=True
    close[oven_141,kitchen_counter_129]=True
    close[oven_141,cupboard_130]=True
    close[oven_141,cupboard_131]=True
    close[oven_141,kitchen_counter_132]=True
    close[oven_141,faucet_134]=True
    close[oven_141,stovefan_139]=True
    close[dishwasher_143,wall_7]=True
    close[dishwasher_143,wall_8]=True
    close[dishwasher_143,floor_21]=True
    close[dishwasher_143,floor_22]=True
    close[dishwasher_143,walllamp_44]=True
    close[dishwasher_143,kitchen_counter_129]=True
    close[dishwasher_143,cupboard_131]=True
    close[dishwasher_143,toaster_144]=True
    close[dishwasher_143,coffe_maker_147]=True
    close[toaster_144,wall_7]=True
    close[toaster_144,wall_8]=True
    close[toaster_144,floor_21]=True
    close[toaster_144,floor_22]=True
    close[toaster_144,ceiling_33]=True
    close[toaster_144,ceiling_34]=True
    close[toaster_144,walllamp_44]=True
    close[toaster_144,kitchen_counter_129]=True
    close[toaster_144,cupboard_131]=True
    close[toaster_144,fridge_140]=True
    close[toaster_144,dishwasher_143]=True
    close[toaster_144,coffe_maker_147]=True
    close[coffe_maker_147,wall_7]=True
    close[coffe_maker_147,wall_8]=True
    close[coffe_maker_147,floor_21]=True
    close[coffe_maker_147,ceiling_33]=True
    close[coffe_maker_147,ceiling_34]=True
    close[coffe_maker_147,walllamp_44]=True
    close[coffe_maker_147,kitchen_counter_129]=True
    close[coffe_maker_147,cupboard_131]=True
    close[coffe_maker_147,dishwasher_143]=True
    close[coffe_maker_147,toaster_144]=True
    close[microwave_149,wall_2]=True
    close[microwave_149,wall_6]=True
    close[microwave_149,floor_15]=True
    close[microwave_149,ceiling_27]=True
    close[microwave_149,walllamp_45]=True
    close[microwave_149,kitchen_counter_128]=True
    close[microwave_149,cupboard_130]=True
    close[microwave_149,kitchen_counter_132]=True
    close[microwave_149,sink_133]=True
    close[microwave_149,faucet_134]=True
    close[microwave_149,wall_172]=True
    close[floor_162,floor_163]=True
    close[floor_162,floor_166]=True
    close[floor_162,floor_168]=True
    close[floor_162,wall_169]=True
    close[floor_162,wall_171]=True
    close[floor_162,tvstand_186]=True
    close[floor_162,wallshelf_187]=True
    close[floor_162,wallshelf_190]=True
    close[floor_162,photoframe_210]=True
    close[floor_162,television_216]=True
    close[floor_162,wall_267]=True
    close[floor_162,floor_278]=True
    close[floor_162,walllamp_291]=True
    close[floor_162,shower_303]=True
    close[floor_162,curtain_304]=True
    close[floor_163,floor_162]=True
    close[floor_163,floor_166]=True
    close[floor_163,floor_168]=True
    close[floor_163,wall_169]=True
    close[floor_163,wall_171]=True
    close[floor_163,tvstand_186]=True
    close[floor_163,wallshelf_187]=True
    close[floor_163,wallshelf_190]=True
    close[floor_163,photoframe_210]=True
    close[floor_163,television_216]=True
    close[floor_163,wall_267]=True
    close[floor_163,floor_278]=True
    close[floor_163,walllamp_291]=True
    close[floor_163,shower_303]=True
    close[floor_163,curtain_304]=True
    close[floor_164,floor_165]=True
    close[floor_164,floor_168]=True
    close[floor_164,wall_170]=True
    close[floor_164,wall_174]=True
    close[floor_164,couch_192]=True
    close[floor_164,table_193]=True
    close[floor_164,orchid_200]=True
    close[floor_164,door_234]=True
    close[floor_164,light_258]=True
    close[floor_165,kitchen_counter_128]=True
    close[floor_165,floor_164]=True
    close[floor_165,floor_167]=True
    close[floor_165,wall_170]=True
    close[floor_165,wall_174]=True
    close[floor_165,doorjamb_182]=True
    close[floor_165,bookshelf_188]=True
    close[floor_165,couch_192]=True
    close[floor_165,table_193]=True
    close[floor_165,orchid_200]=True
    close[floor_165,floor_224]=True
    close[floor_165,wall_232]=True
    close[floor_165,door_234]=True
    close[floor_165,light_258]=True
    close[floor_165,desk_261]=True
    close[floor_166,wall_3]=True
    close[floor_166,floor_14]=True
    close[floor_166,doorjamb_37]=True
    close[floor_166,powersocket_48]=True
    close[floor_166,light_49]=True
    close[floor_166,floor_162]=True
    close[floor_166,floor_163]=True
    close[floor_166,floor_167]=True
    close[floor_166,wall_169]=True
    close[floor_166,wall_171]=True
    close[floor_166,tvstand_186]=True
    close[floor_166,bookshelf_189]=True
    close[floor_166,television_216]=True
    close[floor_166,light_217]=True
    close[floor_166,powersocket_218]=True
    close[floor_166,wall_268]=True
    close[floor_166,floor_277]=True
    close[floor_166,walllamp_291]=True
    close[floor_166,toilet_302]=True
    close[floor_167,wall_6]=True
    close[floor_167,floor_15]=True
    close[floor_167,kitchen_counter_128]=True
    close[floor_167,floor_165]=True
    close[floor_167,floor_166]=True
    close[floor_167,floor_168]=True
    close[floor_167,wall_171]=True
    close[floor_167,wall_172]=True
    close[floor_167,wall_174]=True
    close[floor_167,bookshelf_188]=True
    close[floor_167,bookshelf_189]=True
    close[floor_167,table_193]=True
    close[floor_167,orchid_200]=True
    close[floor_167,light_217]=True
    close[floor_167,powersocket_218]=True
    close[floor_168,floor_162]=True
    close[floor_168,floor_163]=True
    close[floor_168,floor_164]=True
    close[floor_168,floor_167]=True
    close[floor_168,wall_169]=True
    close[floor_168,wall_170]=True
    close[floor_168,wall_173]=True
    close[floor_168,window_181]=True
    close[floor_168,wallshelf_187]=True
    close[floor_168,table_193]=True
    close[floor_168,curtain_197]=True
    close[floor_168,curtain_198]=True
    close[floor_168,curtain_199]=True
    close[floor_168,orchid_200]=True
    close[floor_168,photoframe_210]=True
    close[wall_169,floor_162]=True
    close[wall_169,floor_163]=True
    close[wall_169,floor_166]=True
    close[wall_169,floor_168]=True
    close[wall_169,wall_171]=True
    close[wall_169,wall_173]=True
    close[wall_169,ceiling_175]=True
    close[wall_169,ceiling_176]=True
    close[wall_169,ceiling_178]=True
    close[wall_169,window_181]=True
    close[wall_169,walllamp_184]=True
    close[wall_169,tvstand_186]=True
    close[wall_169,wallshelf_187]=True
    close[wall_169,wallshelf_190]=True
    close[wall_169,wallshelf_191]=True
    close[wall_169,curtain_197]=True
    close[wall_169,curtain_198]=True
    close[wall_169,photoframe_210]=True
    close[wall_169,television_216]=True
    close[wall_169,wall_267]=True
    close[wall_169,floor_278]=True
    close[wall_169,ceiling_282]=True
    close[wall_169,walllamp_291]=True
    close[wall_169,shower_303]=True
    close[wall_169,curtain_304]=True
    close[wall_170,floor_164]=True
    close[wall_170,floor_165]=True
    close[wall_170,floor_168]=True
    close[wall_170,wall_173]=True
    close[wall_170,wall_174]=True
    close[wall_170,ceiling_178]=True
    close[wall_170,ceiling_179]=True
    close[wall_170,ceiling_180]=True
    close[wall_170,window_181]=True
    close[wall_170,doorjamb_182]=True
    close[wall_170,ceilinglamp_185]=True
    close[wall_170,couch_192]=True
    close[wall_170,table_193]=True
    close[wall_170,curtain_199]=True
    close[wall_170,orchid_200]=True
    close[wall_170,door_234]=True
    close[wall_170,light_258]=True
    close[wall_171,wall_3]=True
    close[wall_171,floor_14]=True
    close[wall_171,ceiling_26]=True
    close[wall_171,doorjamb_37]=True
    close[wall_171,powersocket_48]=True
    close[wall_171,light_49]=True
    close[wall_171,floor_162]=True
    close[wall_171,floor_163]=True
    close[wall_171,floor_166]=True
    close[wall_171,floor_167]=True
    close[wall_171,wall_169]=True
    close[wall_171,wall_172]=True
    close[wall_171,ceiling_175]=True
    close[wall_171,ceiling_176]=True
    close[wall_171,ceiling_177]=True
    close[wall_171,walllamp_183]=True
    close[wall_171,tvstand_186]=True
    close[wall_171,bookshelf_189]=True
    close[wall_171,television_216]=True
    close[wall_171,light_217]=True
    close[wall_171,powersocket_218]=True
    close[wall_171,wall_268]=True
    close[wall_171,floor_277]=True
    close[wall_171,ceiling_281]=True
    close[wall_171,walllamp_291]=True
    close[wall_171,toilet_302]=True
    close[wall_171,curtain_304]=True
    close[wall_172,wall_3]=True
    close[wall_172,wall_6]=True
    close[wall_172,floor_15]=True
    close[wall_172,ceiling_27]=True
    close[wall_172,doorjamb_37]=True
    close[wall_172,kitchen_counter_128]=True
    close[wall_172,cupboard_130]=True
    close[wall_172,kitchen_counter_132]=True
    close[wall_172,microwave_149]=True
    close[wall_172,floor_167]=True
    close[wall_172,wall_171]=True
    close[wall_172,wall_174]=True
    close[wall_172,ceiling_177]=True
    close[wall_172,bookshelf_188]=True
    close[wall_172,bookshelf_189]=True
    close[wall_172,light_217]=True
    close[wall_172,powersocket_218]=True
    close[wall_173,floor_168]=True
    close[wall_173,wall_169]=True
    close[wall_173,wall_170]=True
    close[wall_173,ceiling_178]=True
    close[wall_173,window_181]=True
    close[wall_173,wallshelf_187]=True
    close[wall_173,wallshelf_190]=True
    close[wall_173,wallshelf_191]=True
    close[wall_173,curtain_197]=True
    close[wall_173,curtain_198]=True
    close[wall_173,curtain_199]=True
    close[wall_173,photoframe_210]=True
    close[wall_174,kitchen_counter_128]=True
    close[wall_174,floor_164]=True
    close[wall_174,floor_165]=True
    close[wall_174,floor_167]=True
    close[wall_174,wall_170]=True
    close[wall_174,wall_172]=True
    close[wall_174,ceiling_177]=True
    close[wall_174,ceiling_179]=True
    close[wall_174,ceiling_180]=True
    close[wall_174,doorjamb_182]=True
    close[wall_174,ceilinglamp_185]=True
    close[wall_174,bookshelf_188]=True
    close[wall_174,couch_192]=True
    close[wall_174,table_193]=True
    close[wall_174,orchid_200]=True
    close[wall_174,floor_224]=True
    close[wall_174,ceiling_228]=True
    close[wall_174,wall_232]=True
    close[wall_174,door_234]=True
    close[wall_174,light_258]=True
    close[wall_174,desk_261]=True
    close[ceiling_175,wall_169]=True
    close[ceiling_175,wall_171]=True
    close[ceiling_175,ceiling_176]=True
    close[ceiling_175,ceiling_178]=True
    close[ceiling_175,walllamp_184]=True
    close[ceiling_175,wallshelf_190]=True
    close[ceiling_175,wallshelf_191]=True
    close[ceiling_175,curtain_197]=True
    close[ceiling_175,curtain_198]=True
    close[ceiling_175,television_216]=True
    close[ceiling_175,wall_267]=True
    close[ceiling_175,ceiling_282]=True
    close[ceiling_175,walllamp_291]=True
    close[ceiling_175,shower_303]=True
    close[ceiling_175,curtain_304]=True
    close[ceiling_176,wall_3]=True
    close[ceiling_176,ceiling_26]=True
    close[ceiling_176,doorjamb_37]=True
    close[ceiling_176,light_49]=True
    close[ceiling_176,wall_169]=True
    close[ceiling_176,wall_171]=True
    close[ceiling_176,ceiling_175]=True
    close[ceiling_176,ceiling_177]=True
    close[ceiling_176,walllamp_183]=True
    close[ceiling_176,bookshelf_189]=True
    close[ceiling_176,television_216]=True
    close[ceiling_176,light_217]=True
    close[ceiling_176,wall_268]=True
    close[ceiling_176,ceiling_281]=True
    close[ceiling_176,walllamp_291]=True
    close[ceiling_177,wall_6]=True
    close[ceiling_177,ceiling_27]=True
    close[ceiling_177,wall_171]=True
    close[ceiling_177,wall_172]=True
    close[ceiling_177,wall_174]=True
    close[ceiling_177,ceiling_176]=True
    close[ceiling_177,ceiling_178]=True
    close[ceiling_177,ceiling_180]=True
    close[ceiling_177,ceilinglamp_185]=True
    close[ceiling_177,bookshelf_188]=True
    close[ceiling_177,bookshelf_189]=True
    close[ceiling_177,light_217]=True
    close[ceiling_178,wall_169]=True
    close[ceiling_178,wall_170]=True
    close[ceiling_178,wall_173]=True
    close[ceiling_178,ceiling_175]=True
    close[ceiling_178,ceiling_177]=True
    close[ceiling_178,ceiling_179]=True
    close[ceiling_178,window_181]=True
    close[ceiling_178,ceilinglamp_185]=True
    close[ceiling_178,curtain_197]=True
    close[ceiling_178,curtain_198]=True
    close[ceiling_178,curtain_199]=True
    close[ceiling_179,wall_170]=True
    close[ceiling_179,wall_174]=True
    close[ceiling_179,ceiling_178]=True
    close[ceiling_179,ceiling_180]=True
    close[ceiling_179,ceilinglamp_185]=True
    close[ceiling_179,couch_192]=True
    close[ceiling_179,curtain_199]=True
    close[ceiling_179,light_258]=True
    close[ceiling_180,wall_170]=True
    close[ceiling_180,wall_174]=True
    close[ceiling_180,ceiling_177]=True
    close[ceiling_180,ceiling_179]=True
    close[ceiling_180,doorjamb_182]=True
    close[ceiling_180,ceilinglamp_185]=True
    close[ceiling_180,bookshelf_188]=True
    close[ceiling_180,ceiling_228]=True
    close[ceiling_180,wall_232]=True
    close[ceiling_180,light_258]=True
    close[window_181,floor_168]=True
    close[window_181,wall_169]=True
    close[window_181,wall_170]=True
    close[window_181,wall_173]=True
    close[window_181,ceiling_178]=True
    close[window_181,wallshelf_187]=True
    close[window_181,wallshelf_190]=True
    close[window_181,wallshelf_191]=True
    close[window_181,curtain_197]=True
    close[window_181,curtain_198]=True
    close[window_181,curtain_199]=True
    close[window_181,photoframe_210]=True
    close[doorjamb_182,floor_165]=True
    close[doorjamb_182,wall_170]=True
    close[doorjamb_182,wall_174]=True
    close[doorjamb_182,ceiling_180]=True
    close[doorjamb_182,bookshelf_188]=True
    close[doorjamb_182,couch_192]=True
    close[doorjamb_182,floor_224]=True
    close[doorjamb_182,ceiling_228]=True
    close[doorjamb_182,wall_231]=True
    close[doorjamb_182,wall_232]=True
    close[doorjamb_182,door_234]=True
    close[doorjamb_182,light_258]=True
    close[doorjamb_182,desk_261]=True
    close[walllamp_183,wall_3]=True
    close[walllamp_183,wall_5]=True
    close[walllamp_183,ceiling_25]=True
    close[walllamp_183,ceiling_26]=True
    close[walllamp_183,doorjamb_37]=True
    close[walllamp_183,light_49]=True
    close[walllamp_183,wall_171]=True
    close[walllamp_183,ceiling_176]=True
    close[walllamp_183,tvstand_186]=True
    close[walllamp_183,television_216]=True
    close[walllamp_183,wall_268]=True
    close[walllamp_183,ceiling_281]=True
    close[walllamp_183,walllamp_291]=True
    close[walllamp_183,toilet_302]=True
    close[walllamp_184,wall_169]=True
    close[walllamp_184,ceiling_175]=True
    close[walllamp_184,tvstand_186]=True
    close[walllamp_184,wallshelf_187]=True
    close[walllamp_184,wallshelf_190]=True
    close[walllamp_184,wallshelf_191]=True
    close[walllamp_184,television_216]=True
    close[walllamp_184,wall_267]=True
    close[walllamp_184,ceiling_282]=True
    close[walllamp_184,walllamp_291]=True
    close[walllamp_184,shower_303]=True
    close[walllamp_184,curtain_304]=True
    close[ceilinglamp_185,wall_170]=True
    close[ceilinglamp_185,wall_174]=True
    close[ceilinglamp_185,ceiling_177]=True
    close[ceilinglamp_185,ceiling_178]=True
    close[ceilinglamp_185,ceiling_179]=True
    close[ceilinglamp_185,ceiling_180]=True
    close[tvstand_186,powersocket_48]=True
    close[tvstand_186,floor_162]=True
    close[tvstand_186,floor_163]=True
    close[tvstand_186,floor_166]=True
    close[tvstand_186,wall_169]=True
    close[tvstand_186,wall_171]=True
    close[tvstand_186,walllamp_183]=True
    close[tvstand_186,walllamp_184]=True
    close[tvstand_186,wallshelf_187]=True
    close[tvstand_186,wallshelf_190]=True
    close[tvstand_186,photoframe_210]=True
    close[tvstand_186,television_216]=True
    close[tvstand_186,wall_267]=True
    close[tvstand_186,wall_268]=True
    close[tvstand_186,floor_277]=True
    close[tvstand_186,floor_278]=True
    close[tvstand_186,walllamp_291]=True
    close[tvstand_186,toilet_302]=True
    close[tvstand_186,shower_303]=True
    close[tvstand_186,curtain_304]=True
    close[wallshelf_187,floor_162]=True
    close[wallshelf_187,floor_163]=True
    close[wallshelf_187,floor_168]=True
    close[wallshelf_187,wall_169]=True
    close[wallshelf_187,wall_173]=True
    close[wallshelf_187,window_181]=True
    close[wallshelf_187,walllamp_184]=True
    close[wallshelf_187,tvstand_186]=True
    close[wallshelf_187,wallshelf_190]=True
    close[wallshelf_187,wallshelf_191]=True
    close[wallshelf_187,curtain_197]=True
    close[wallshelf_187,curtain_198]=True
    close[wallshelf_187,photoframe_210]=True
    close[wallshelf_187,wall_267]=True
    close[wallshelf_187,floor_278]=True
    close[wallshelf_187,shower_303]=True
    close[bookshelf_188,wall_6]=True
    close[bookshelf_188,floor_15]=True
    close[bookshelf_188,kitchen_counter_128]=True
    close[bookshelf_188,floor_165]=True
    close[bookshelf_188,floor_167]=True
    close[bookshelf_188,wall_172]=True
    close[bookshelf_188,wall_174]=True
    close[bookshelf_188,ceiling_177]=True
    close[bookshelf_188,ceiling_180]=True
    close[bookshelf_188,doorjamb_182]=True
    close[bookshelf_188,bookshelf_189]=True
    close[bookshelf_188,door_234]=True
    close[bookshelf_189,wall_3]=True
    close[bookshelf_189,wall_6]=True
    close[bookshelf_189,floor_14]=True
    close[bookshelf_189,floor_15]=True
    close[bookshelf_189,ceiling_27]=True
    close[bookshelf_189,doorjamb_37]=True
    close[bookshelf_189,kitchen_counter_128]=True
    close[bookshelf_189,floor_166]=True
    close[bookshelf_189,floor_167]=True
    close[bookshelf_189,wall_171]=True
    close[bookshelf_189,wall_172]=True
    close[bookshelf_189,ceiling_176]=True
    close[bookshelf_189,ceiling_177]=True
    close[bookshelf_189,bookshelf_188]=True
    close[bookshelf_189,light_217]=True
    close[bookshelf_189,powersocket_218]=True
    close[wallshelf_190,floor_162]=True
    close[wallshelf_190,floor_163]=True
    close[wallshelf_190,wall_169]=True
    close[wallshelf_190,wall_173]=True
    close[wallshelf_190,ceiling_175]=True
    close[wallshelf_190,window_181]=True
    close[wallshelf_190,walllamp_184]=True
    close[wallshelf_190,tvstand_186]=True
    close[wallshelf_190,wallshelf_187]=True
    close[wallshelf_190,wallshelf_191]=True
    close[wallshelf_190,curtain_197]=True
    close[wallshelf_190,curtain_198]=True
    close[wallshelf_190,photoframe_210]=True
    close[wallshelf_190,wall_267]=True
    close[wallshelf_190,shower_303]=True
    close[wallshelf_191,wall_169]=True
    close[wallshelf_191,wall_173]=True
    close[wallshelf_191,ceiling_175]=True
    close[wallshelf_191,window_181]=True
    close[wallshelf_191,walllamp_184]=True
    close[wallshelf_191,wallshelf_187]=True
    close[wallshelf_191,wallshelf_190]=True
    close[wallshelf_191,curtain_197]=True
    close[wallshelf_191,curtain_198]=True
    close[wallshelf_191,photoframe_210]=True
    close[wallshelf_191,wall_267]=True
    close[wallshelf_191,shower_303]=True
    close[couch_192,floor_164]=True
    close[couch_192,floor_165]=True
    close[couch_192,wall_170]=True
    close[couch_192,wall_174]=True
    close[couch_192,ceiling_179]=True
    close[couch_192,doorjamb_182]=True
    close[couch_192,table_193]=True
    close[couch_192,orchid_200]=True
    close[couch_192,television_216]=True
    close[couch_192,floor_224]=True
    close[couch_192,wall_232]=True
    close[couch_192,door_234]=True
    close[couch_192,light_258]=True
    close[table_193,computer_2110]=True
    close[table_193,floor_164]=True
    close[table_193,floor_165]=True
    close[table_193,floor_167]=True
    close[table_193,floor_168]=True
    close[table_193,wall_170]=True
    close[table_193,wall_174]=True
    close[table_193,couch_192]=True
    close[table_193,curtain_199]=True
    close[table_193,orchid_200]=True
    close[curtain_197,floor_168]=True
    close[curtain_197,wall_169]=True
    close[curtain_197,wall_173]=True
    close[curtain_197,ceiling_175]=True
    close[curtain_197,ceiling_178]=True
    close[curtain_197,window_181]=True
    close[curtain_197,wallshelf_187]=True
    close[curtain_197,wallshelf_190]=True
    close[curtain_197,wallshelf_191]=True
    close[curtain_197,curtain_198]=True
    close[curtain_197,curtain_199]=True
    close[curtain_197,photoframe_210]=True
    close[curtain_198,floor_168]=True
    close[curtain_198,wall_169]=True
    close[curtain_198,wall_173]=True
    close[curtain_198,ceiling_175]=True
    close[curtain_198,ceiling_178]=True
    close[curtain_198,window_181]=True
    close[curtain_198,wallshelf_187]=True
    close[curtain_198,wallshelf_190]=True
    close[curtain_198,wallshelf_191]=True
    close[curtain_198,curtain_197]=True
    close[curtain_198,curtain_199]=True
    close[curtain_198,photoframe_210]=True
    close[curtain_199,floor_168]=True
    close[curtain_199,wall_170]=True
    close[curtain_199,wall_173]=True
    close[curtain_199,ceiling_178]=True
    close[curtain_199,ceiling_179]=True
    close[curtain_199,window_181]=True
    close[curtain_199,table_193]=True
    close[curtain_199,curtain_197]=True
    close[curtain_199,curtain_198]=True
    close[orchid_200,floor_164]=True
    close[orchid_200,floor_165]=True
    close[orchid_200,floor_167]=True
    close[orchid_200,floor_168]=True
    close[orchid_200,wall_170]=True
    close[orchid_200,wall_174]=True
    close[orchid_200,couch_192]=True
    close[orchid_200,table_193]=True
    close[photoframe_210,floor_162]=True
    close[photoframe_210,floor_163]=True
    close[photoframe_210,floor_168]=True
    close[photoframe_210,wall_169]=True
    close[photoframe_210,wall_173]=True
    close[photoframe_210,window_181]=True
    close[photoframe_210,tvstand_186]=True
    close[photoframe_210,wallshelf_187]=True
    close[photoframe_210,wallshelf_190]=True
    close[photoframe_210,wallshelf_191]=True
    close[photoframe_210,curtain_197]=True
    close[photoframe_210,curtain_198]=True
    close[television_216,floor_162]=True
    close[television_216,floor_163]=True
    close[television_216,floor_166]=True
    close[television_216,wall_169]=True
    close[television_216,wall_171]=True
    close[television_216,ceiling_175]=True
    close[television_216,ceiling_176]=True
    close[television_216,walllamp_183]=True
    close[television_216,walllamp_184]=True
    close[television_216,tvstand_186]=True
    close[television_216,couch_192]=True
    close[television_216,wall_267]=True
    close[television_216,wall_268]=True
    close[television_216,floor_277]=True
    close[television_216,floor_278]=True
    close[television_216,walllamp_291]=True
    close[television_216,shower_303]=True
    close[television_216,curtain_304]=True
    close[light_217,wall_3]=True
    close[light_217,wall_6]=True
    close[light_217,floor_14]=True
    close[light_217,floor_15]=True
    close[light_217,ceiling_26]=True
    close[light_217,ceiling_27]=True
    close[light_217,doorjamb_37]=True
    close[light_217,powersocket_48]=True
    close[light_217,light_49]=True
    close[light_217,floor_166]=True
    close[light_217,floor_167]=True
    close[light_217,wall_171]=True
    close[light_217,wall_172]=True
    close[light_217,ceiling_176]=True
    close[light_217,ceiling_177]=True
    close[light_217,bookshelf_189]=True
    close[light_217,powersocket_218]=True
    close[powersocket_218,wall_3]=True
    close[powersocket_218,wall_6]=True
    close[powersocket_218,floor_14]=True
    close[powersocket_218,floor_15]=True
    close[powersocket_218,doorjamb_37]=True
    close[powersocket_218,powersocket_48]=True
    close[powersocket_218,light_49]=True
    close[powersocket_218,floor_166]=True
    close[powersocket_218,floor_167]=True
    close[powersocket_218,wall_171]=True
    close[powersocket_218,wall_172]=True
    close[powersocket_218,bookshelf_189]=True
    close[powersocket_218,light_217]=True
    close[bedroom_220,ironing_board_2099]=True
    close[floor_221,floor_222]=True
    close[floor_221,floor_223]=True
    close[floor_221,floor_225]=True
    close[floor_221,wall_230]=True
    close[floor_221,wall_231]=True
    close[floor_221,wall_233]=True
    close[floor_221,tablelamp_236]=True
    close[floor_221,photoframe_246]=True
    close[floor_221,powersocket_259]=True
    close[floor_221,bookshelf_260]=True
    close[floor_221,nightstand_262]=True
    close[floor_221,bed_264]=True
    close[floor_222,floor_221]=True
    close[floor_222,floor_223]=True
    close[floor_222,floor_225]=True
    close[floor_222,wall_230]=True
    close[floor_222,wall_231]=True
    close[floor_222,wall_233]=True
    close[floor_222,tablelamp_236]=True
    close[floor_222,photoframe_246]=True
    close[floor_222,powersocket_259]=True
    close[floor_222,bookshelf_260]=True
    close[floor_222,nightstand_262]=True
    close[floor_222,bed_264]=True
    close[floor_223,floor_221]=True
    close[floor_223,floor_222]=True
    close[floor_223,floor_224]=True
    close[floor_223,wall_231]=True
    close[floor_223,wall_232]=True
    close[floor_223,wall_233]=True
    close[floor_223,door_234]=True
    close[floor_223,photoframe_246]=True
    close[floor_223,bookshelf_260]=True
    close[floor_223,desk_261]=True
    close[floor_224,floor_165]=True
    close[floor_224,wall_174]=True
    close[floor_224,doorjamb_182]=True
    close[floor_224,couch_192]=True
    close[floor_224,floor_223]=True
    close[floor_224,floor_225]=True
    close[floor_224,wall_230]=True
    close[floor_224,wall_231]=True
    close[floor_224,wall_232]=True
    close[floor_224,door_234]=True
    close[floor_224,light_258]=True
    close[floor_224,desk_261]=True
    close[floor_224,bed_264]=True
    close[floor_225,floor_221]=True
    close[floor_225,floor_222]=True
    close[floor_225,floor_224]=True
    close[floor_225,wall_230]=True
    close[floor_225,wall_232]=True
    close[floor_225,wall_233]=True
    close[floor_225,tablelamp_236]=True
    close[floor_225,nightstand_262]=True
    close[floor_225,bed_264]=True
    close[ceiling_226,ceiling_227]=True
    close[ceiling_226,ceiling_229]=True
    close[ceiling_226,wall_230]=True
    close[ceiling_226,wall_231]=True
    close[ceiling_226,wall_233]=True
    close[ceiling_226,ceilinglamp_235]=True
    close[ceiling_226,photoframe_246]=True
    close[ceiling_226,bookshelf_260]=True
    close[ceiling_227,ceiling_226]=True
    close[ceiling_227,ceiling_228]=True
    close[ceiling_227,wall_231]=True
    close[ceiling_227,wall_232]=True
    close[ceiling_227,wall_233]=True
    close[ceiling_227,ceilinglamp_235]=True
    close[ceiling_227,photoframe_246]=True
    close[ceiling_227,bookshelf_260]=True
    close[ceiling_228,wall_174]=True
    close[ceiling_228,ceiling_180]=True
    close[ceiling_228,doorjamb_182]=True
    close[ceiling_228,ceiling_227]=True
    close[ceiling_228,ceiling_229]=True
    close[ceiling_228,wall_230]=True
    close[ceiling_228,wall_231]=True
    close[ceiling_228,wall_232]=True
    close[ceiling_228,ceilinglamp_235]=True
    close[ceiling_228,light_258]=True
    close[ceiling_229,ceiling_226]=True
    close[ceiling_229,ceiling_228]=True
    close[ceiling_229,wall_230]=True
    close[ceiling_229,wall_232]=True
    close[ceiling_229,wall_233]=True
    close[ceiling_229,ceilinglamp_235]=True
    close[wall_230,floor_221]=True
    close[wall_230,floor_222]=True
    close[wall_230,floor_224]=True
    close[wall_230,floor_225]=True
    close[wall_230,ceiling_226]=True
    close[wall_230,ceiling_228]=True
    close[wall_230,ceiling_229]=True
    close[wall_230,wall_232]=True
    close[wall_230,wall_233]=True
    close[wall_230,ceilinglamp_235]=True
    close[wall_230,tablelamp_236]=True
    close[wall_230,nightstand_262]=True
    close[wall_230,bed_264]=True
    close[wall_231,doorjamb_182]=True
    close[wall_231,floor_221]=True
    close[wall_231,floor_222]=True
    close[wall_231,floor_223]=True
    close[wall_231,floor_224]=True
    close[wall_231,ceiling_226]=True
    close[wall_231,ceiling_227]=True
    close[wall_231,ceiling_228]=True
    close[wall_231,wall_232]=True
    close[wall_231,wall_233]=True
    close[wall_231,door_234]=True
    close[wall_231,ceilinglamp_235]=True
    close[wall_231,photoframe_246]=True
    close[wall_231,bookshelf_260]=True
    close[wall_231,desk_261]=True
    close[wall_232,floor_165]=True
    close[wall_232,wall_174]=True
    close[wall_232,ceiling_180]=True
    close[wall_232,doorjamb_182]=True
    close[wall_232,couch_192]=True
    close[wall_232,floor_223]=True
    close[wall_232,floor_224]=True
    close[wall_232,floor_225]=True
    close[wall_232,ceiling_227]=True
    close[wall_232,ceiling_228]=True
    close[wall_232,ceiling_229]=True
    close[wall_232,wall_230]=True
    close[wall_232,wall_231]=True
    close[wall_232,door_234]=True
    close[wall_232,ceilinglamp_235]=True
    close[wall_232,light_258]=True
    close[wall_232,desk_261]=True
    close[wall_232,bed_264]=True
    close[wall_233,floor_221]=True
    close[wall_233,floor_222]=True
    close[wall_233,floor_223]=True
    close[wall_233,floor_225]=True
    close[wall_233,ceiling_226]=True
    close[wall_233,ceiling_227]=True
    close[wall_233,ceiling_229]=True
    close[wall_233,wall_230]=True
    close[wall_233,wall_231]=True
    close[wall_233,ceilinglamp_235]=True
    close[wall_233,tablelamp_236]=True
    close[wall_233,photoframe_246]=True
    close[wall_233,powersocket_259]=True
    close[wall_233,bookshelf_260]=True
    close[wall_233,nightstand_262]=True
    close[wall_233,bed_264]=True
    close[door_234,floor_164]=True
    close[door_234,floor_165]=True
    close[door_234,wall_170]=True
    close[door_234,wall_174]=True
    close[door_234,doorjamb_182]=True
    close[door_234,bookshelf_188]=True
    close[door_234,couch_192]=True
    close[door_234,floor_223]=True
    close[door_234,floor_224]=True
    close[door_234,wall_231]=True
    close[door_234,wall_232]=True
    close[door_234,light_258]=True
    close[door_234,desk_261]=True
    close[ceilinglamp_235,ceiling_226]=True
    close[ceilinglamp_235,ceiling_227]=True
    close[ceilinglamp_235,ceiling_228]=True
    close[ceilinglamp_235,ceiling_229]=True
    close[ceilinglamp_235,wall_230]=True
    close[ceilinglamp_235,wall_231]=True
    close[ceilinglamp_235,wall_232]=True
    close[ceilinglamp_235,wall_233]=True
    close[tablelamp_236,floor_221]=True
    close[tablelamp_236,floor_222]=True
    close[tablelamp_236,floor_225]=True
    close[tablelamp_236,wall_230]=True
    close[tablelamp_236,wall_233]=True
    close[tablelamp_236,nightstand_262]=True
    close[tablelamp_236,bed_264]=True
    close[photoframe_246,floor_221]=True
    close[photoframe_246,floor_222]=True
    close[photoframe_246,floor_223]=True
    close[photoframe_246,ceiling_226]=True
    close[photoframe_246,ceiling_227]=True
    close[photoframe_246,wall_231]=True
    close[photoframe_246,wall_233]=True
    close[photoframe_246,bookshelf_260]=True
    close[photoframe_246,desk_261]=True
    close[light_258,floor_164]=True
    close[light_258,floor_165]=True
    close[light_258,wall_170]=True
    close[light_258,wall_174]=True
    close[light_258,ceiling_179]=True
    close[light_258,ceiling_180]=True
    close[light_258,doorjamb_182]=True
    close[light_258,couch_192]=True
    close[light_258,floor_224]=True
    close[light_258,ceiling_228]=True
    close[light_258,wall_232]=True
    close[light_258,door_234]=True
    close[powersocket_259,floor_221]=True
    close[powersocket_259,floor_222]=True
    close[powersocket_259,wall_233]=True
    close[powersocket_259,bookshelf_260]=True
    close[powersocket_259,nightstand_262]=True
    close[bookshelf_260,floor_221]=True
    close[bookshelf_260,floor_222]=True
    close[bookshelf_260,floor_223]=True
    close[bookshelf_260,ceiling_226]=True
    close[bookshelf_260,ceiling_227]=True
    close[bookshelf_260,wall_231]=True
    close[bookshelf_260,wall_233]=True
    close[bookshelf_260,photoframe_246]=True
    close[bookshelf_260,powersocket_259]=True
    close[desk_261,floor_165]=True
    close[desk_261,wall_174]=True
    close[desk_261,doorjamb_182]=True
    close[desk_261,floor_223]=True
    close[desk_261,floor_224]=True
    close[desk_261,wall_231]=True
    close[desk_261,wall_232]=True
    close[desk_261,door_234]=True
    close[desk_261,photoframe_246]=True
    close[nightstand_262,floor_221]=True
    close[nightstand_262,floor_222]=True
    close[nightstand_262,floor_225]=True
    close[nightstand_262,wall_230]=True
    close[nightstand_262,wall_233]=True
    close[nightstand_262,tablelamp_236]=True
    close[nightstand_262,powersocket_259]=True
    close[nightstand_262,bed_264]=True
    close[bed_264,floor_221]=True
    close[bed_264,floor_222]=True
    close[bed_264,floor_224]=True
    close[bed_264,floor_225]=True
    close[bed_264,wall_230]=True
    close[bed_264,wall_232]=True
    close[bed_264,wall_233]=True
    close[bed_264,tablelamp_236]=True
    close[bed_264,nightstand_262]=True
    close[wall_266,wall_269]=True
    close[wall_266,wall_270]=True
    close[wall_266,floor_272]=True
    close[wall_266,floor_273]=True
    close[wall_266,floor_274]=True
    close[wall_266,floor_275]=True
    close[wall_266,ceiling_279]=True
    close[wall_266,ceiling_283]=True
    close[wall_266,ceiling_284]=True
    close[wall_266,window_287]=True
    close[wall_266,ceilinglamp_288]=True
    close[wall_266,walllamp_289]=True
    close[wall_266,bathtub_297]=True
    close[wall_266,wallshelf_301]=True
    close[wall_266,bathroom_cabinet_305]=True
    close[wall_266,bathroom_counter_306]=True
    close[wall_266,sink_307]=True
    close[wall_266,faucet_308]=True
    close[wall_267,floor_162]=True
    close[wall_267,floor_163]=True
    close[wall_267,wall_169]=True
    close[wall_267,ceiling_175]=True
    close[wall_267,walllamp_184]=True
    close[wall_267,tvstand_186]=True
    close[wall_267,wallshelf_187]=True
    close[wall_267,wallshelf_190]=True
    close[wall_267,wallshelf_191]=True
    close[wall_267,television_216]=True
    close[wall_267,wall_268]=True
    close[wall_267,wall_270]=True
    close[wall_267,floor_275]=True
    close[wall_267,floor_277]=True
    close[wall_267,floor_278]=True
    close[wall_267,ceiling_281]=True
    close[wall_267,ceiling_282]=True
    close[wall_267,ceiling_283]=True
    close[wall_267,window_287]=True
    close[wall_267,ceilinglamp_288]=True
    close[wall_267,walllamp_291]=True
    close[wall_267,curtain_293]=True
    close[wall_267,curtain_294]=True
    close[wall_267,shower_303]=True
    close[wall_267,curtain_304]=True
    close[wall_268,wall_3]=True
    close[wall_268,wall_5]=True
    close[wall_268,floor_12]=True
    close[wall_268,floor_13]=True
    close[wall_268,ceiling_25]=True
    close[wall_268,doorjamb_37]=True
    close[wall_268,powersocket_48]=True
    close[wall_268,light_49]=True
    close[wall_268,floor_166]=True
    close[wall_268,wall_171]=True
    close[wall_268,ceiling_176]=True
    close[wall_268,walllamp_183]=True
    close[wall_268,tvstand_186]=True
    close[wall_268,television_216]=True
    close[wall_268,wall_267]=True
    close[wall_268,wall_271]=True
    close[wall_268,floor_276]=True
    close[wall_268,floor_277]=True
    close[wall_268,floor_278]=True
    close[wall_268,ceiling_280]=True
    close[wall_268,ceiling_281]=True
    close[wall_268,ceiling_282]=True
    close[wall_268,doorjamb_285]=True
    close[wall_268,door_286]=True
    close[wall_268,ceilinglamp_288]=True
    close[wall_268,walllamp_291]=True
    close[wall_268,toilet_302]=True
    close[wall_268,curtain_304]=True
    close[wall_269,wall_266]=True
    close[wall_269,wall_271]=True
    close[wall_269,floor_272]=True
    close[wall_269,floor_273]=True
    close[wall_269,floor_274]=True
    close[wall_269,floor_276]=True
    close[wall_269,ceiling_279]=True
    close[wall_269,ceiling_280]=True
    close[wall_269,ceiling_284]=True
    close[wall_269,doorjamb_285]=True
    close[wall_269,door_286]=True
    close[wall_269,ceilinglamp_288]=True
    close[wall_269,walllamp_290]=True
    close[wall_269,bathroom_cabinet_305]=True
    close[wall_269,bathroom_counter_306]=True
    close[wall_269,sink_307]=True
    close[wall_269,faucet_308]=True
    close[wall_269,light_325]=True
    close[wall_269,floor_332]=True
    close[wall_269,wall_339]=True
    close[wall_269,ceiling_350]=True
    close[wall_269,photoframe_361]=True
    close[wall_269,bookshelf_372]=True
    close[wall_270,wall_266]=True
    close[wall_270,wall_267]=True
    close[wall_270,floor_275]=True
    close[wall_270,ceiling_283]=True
    close[wall_270,window_287]=True
    close[wall_270,curtain_293]=True
    close[wall_270,curtain_294]=True
    close[wall_270,bathtub_297]=True
    close[wall_270,wallshelf_301]=True
    close[wall_271,wall_5]=True
    close[wall_271,wall_268]=True
    close[wall_271,wall_269]=True
    close[wall_271,floor_276]=True
    close[wall_271,ceiling_280]=True
    close[wall_271,doorjamb_285]=True
    close[wall_271,door_286]=True
    close[wall_271,light_325]=True
    close[wall_271,floor_337]=True
    close[wall_271,wall_339]=True
    close[wall_271,wall_345]=True
    close[wall_271,ceiling_355]=True
    close[wall_271,desk_375]=True
    close[floor_272,wall_266]=True
    close[floor_272,wall_269]=True
    close[floor_272,floor_273]=True
    close[floor_272,floor_274]=True
    close[floor_272,floor_276]=True
    close[floor_272,door_286]=True
    close[floor_272,walllamp_290]=True
    close[floor_272,bathroom_counter_306]=True
    close[floor_272,sink_307]=True
    close[floor_272,faucet_308]=True
    close[floor_272,light_325]=True
    close[floor_272,floor_332]=True
    close[floor_272,wall_339]=True
    close[floor_272,bookshelf_372]=True
    close[floor_273,wall_266]=True
    close[floor_273,wall_269]=True
    close[floor_273,floor_272]=True
    close[floor_273,floor_274]=True
    close[floor_273,floor_276]=True
    close[floor_273,door_286]=True
    close[floor_273,walllamp_290]=True
    close[floor_273,bathroom_counter_306]=True
    close[floor_273,sink_307]=True
    close[floor_273,faucet_308]=True
    close[floor_273,light_325]=True
    close[floor_273,floor_332]=True
    close[floor_273,wall_339]=True
    close[floor_273,bookshelf_372]=True
    close[floor_274,wall_266]=True
    close[floor_274,wall_269]=True
    close[floor_274,floor_272]=True
    close[floor_274,floor_273]=True
    close[floor_274,floor_275]=True
    close[floor_274,walllamp_289]=True
    close[floor_274,bathtub_297]=True
    close[floor_274,bathroom_counter_306]=True
    close[floor_274,sink_307]=True
    close[floor_274,faucet_308]=True
    close[floor_275,wall_266]=True
    close[floor_275,wall_267]=True
    close[floor_275,wall_270]=True
    close[floor_275,floor_274]=True
    close[floor_275,floor_276]=True
    close[floor_275,floor_278]=True
    close[floor_275,window_287]=True
    close[floor_275,curtain_293]=True
    close[floor_275,curtain_294]=True
    close[floor_275,bathtub_297]=True
    close[floor_276,wall_268]=True
    close[floor_276,wall_269]=True
    close[floor_276,wall_271]=True
    close[floor_276,floor_272]=True
    close[floor_276,floor_273]=True
    close[floor_276,floor_275]=True
    close[floor_276,floor_277]=True
    close[floor_276,doorjamb_285]=True
    close[floor_276,door_286]=True
    close[floor_276,light_325]=True
    close[floor_276,floor_337]=True
    close[floor_276,wall_345]=True
    close[floor_277,wall_5]=True
    close[floor_277,floor_12]=True
    close[floor_277,floor_13]=True
    close[floor_277,powersocket_48]=True
    close[floor_277,light_49]=True
    close[floor_277,floor_166]=True
    close[floor_277,wall_171]=True
    close[floor_277,tvstand_186]=True
    close[floor_277,television_216]=True
    close[floor_277,wall_267]=True
    close[floor_277,wall_268]=True
    close[floor_277,floor_276]=True
    close[floor_277,floor_278]=True
    close[floor_277,door_286]=True
    close[floor_277,walllamp_291]=True
    close[floor_277,toilet_302]=True
    close[floor_278,floor_162]=True
    close[floor_278,floor_163]=True
    close[floor_278,wall_169]=True
    close[floor_278,tvstand_186]=True
    close[floor_278,wallshelf_187]=True
    close[floor_278,television_216]=True
    close[floor_278,wall_267]=True
    close[floor_278,wall_268]=True
    close[floor_278,floor_275]=True
    close[floor_278,floor_277]=True
    close[floor_278,walllamp_291]=True
    close[floor_278,shower_303]=True
    close[floor_278,curtain_304]=True
    close[ceiling_279,wall_266]=True
    close[ceiling_279,wall_269]=True
    close[ceiling_279,ceiling_280]=True
    close[ceiling_279,ceiling_284]=True
    close[ceiling_279,ceilinglamp_288]=True
    close[ceiling_279,walllamp_290]=True
    close[ceiling_279,bathroom_cabinet_305]=True
    close[ceiling_279,faucet_308]=True
    close[ceiling_279,light_325]=True
    close[ceiling_279,wall_339]=True
    close[ceiling_279,ceiling_350]=True
    close[ceiling_279,photoframe_361]=True
    close[ceiling_279,bookshelf_372]=True
    close[ceiling_280,wall_268]=True
    close[ceiling_280,wall_269]=True
    close[ceiling_280,wall_271]=True
    close[ceiling_280,ceiling_279]=True
    close[ceiling_280,ceiling_281]=True
    close[ceiling_280,ceiling_283]=True
    close[ceiling_280,doorjamb_285]=True
    close[ceiling_280,ceilinglamp_288]=True
    close[ceiling_280,light_325]=True
    close[ceiling_280,wall_345]=True
    close[ceiling_280,ceiling_355]=True
    close[ceiling_281,wall_5]=True
    close[ceiling_281,ceiling_25]=True
    close[ceiling_281,wall_171]=True
    close[ceiling_281,ceiling_176]=True
    close[ceiling_281,walllamp_183]=True
    close[ceiling_281,wall_267]=True
    close[ceiling_281,wall_268]=True
    close[ceiling_281,ceiling_280]=True
    close[ceiling_281,ceiling_282]=True
    close[ceiling_281,ceilinglamp_288]=True
    close[ceiling_281,walllamp_291]=True
    close[ceiling_282,wall_169]=True
    close[ceiling_282,ceiling_175]=True
    close[ceiling_282,walllamp_184]=True
    close[ceiling_282,wall_267]=True
    close[ceiling_282,wall_268]=True
    close[ceiling_282,ceiling_281]=True
    close[ceiling_282,ceiling_283]=True
    close[ceiling_282,ceilinglamp_288]=True
    close[ceiling_282,walllamp_291]=True
    close[ceiling_282,curtain_293]=True
    close[ceiling_282,curtain_294]=True
    close[ceiling_282,shower_303]=True
    close[ceiling_282,curtain_304]=True
    close[ceiling_283,wall_266]=True
    close[ceiling_283,wall_267]=True
    close[ceiling_283,wall_270]=True
    close[ceiling_283,ceiling_280]=True
    close[ceiling_283,ceiling_282]=True
    close[ceiling_283,ceiling_284]=True
    close[ceiling_283,window_287]=True
    close[ceiling_283,ceilinglamp_288]=True
    close[ceiling_283,curtain_293]=True
    close[ceiling_283,curtain_294]=True
    close[ceiling_283,wallshelf_301]=True
    close[ceiling_284,wall_266]=True
    close[ceiling_284,wall_269]=True
    close[ceiling_284,ceiling_279]=True
    close[ceiling_284,ceiling_283]=True
    close[ceiling_284,ceilinglamp_288]=True
    close[ceiling_284,walllamp_289]=True
    close[ceiling_284,wallshelf_301]=True
    close[ceiling_284,bathroom_cabinet_305]=True
    close[doorjamb_285,wall_5]=True
    close[doorjamb_285,bookshelf_136]=True
    close[doorjamb_285,wall_268]=True
    close[doorjamb_285,wall_269]=True
    close[doorjamb_285,wall_271]=True
    close[doorjamb_285,floor_276]=True
    close[doorjamb_285,ceiling_280]=True
    close[doorjamb_285,door_286]=True
    close[doorjamb_285,light_325]=True
    close[doorjamb_285,floor_337]=True
    close[doorjamb_285,wall_339]=True
    close[doorjamb_285,wall_345]=True
    close[doorjamb_285,ceiling_355]=True
    close[doorjamb_285,desk_375]=True
    close[doorjamb_285,computer_379]=True
    close[door_286,wall_5]=True
    close[door_286,floor_12]=True
    close[door_286,floor_13]=True
    close[door_286,bookshelf_136]=True
    close[door_286,wall_268]=True
    close[door_286,wall_269]=True
    close[door_286,wall_271]=True
    close[door_286,floor_272]=True
    close[door_286,floor_273]=True
    close[door_286,floor_276]=True
    close[door_286,floor_277]=True
    close[door_286,doorjamb_285]=True
    close[door_286,light_325]=True
    close[door_286,floor_332]=True
    close[door_286,floor_337]=True
    close[door_286,wall_339]=True
    close[door_286,wall_345]=True
    close[door_286,desk_375]=True
    close[door_286,computer_379]=True
    close[window_287,washing_machine_2041]=True
    close[window_287,wall_266]=True
    close[window_287,wall_267]=True
    close[window_287,wall_270]=True
    close[window_287,floor_275]=True
    close[window_287,ceiling_283]=True
    close[window_287,curtain_293]=True
    close[window_287,curtain_294]=True
    close[window_287,bathtub_297]=True
    close[ceilinglamp_288,wall_266]=True
    close[ceilinglamp_288,wall_267]=True
    close[ceilinglamp_288,wall_268]=True
    close[ceilinglamp_288,wall_269]=True
    close[ceilinglamp_288,ceiling_279]=True
    close[ceilinglamp_288,ceiling_280]=True
    close[ceilinglamp_288,ceiling_281]=True
    close[ceilinglamp_288,ceiling_282]=True
    close[ceilinglamp_288,ceiling_283]=True
    close[ceilinglamp_288,ceiling_284]=True
    close[walllamp_289,wall_266]=True
    close[walllamp_289,floor_274]=True
    close[walllamp_289,ceiling_284]=True
    close[walllamp_289,bathtub_297]=True
    close[walllamp_289,wallshelf_301]=True
    close[walllamp_289,bathroom_cabinet_305]=True
    close[walllamp_289,bathroom_counter_306]=True
    close[walllamp_290,wall_269]=True
    close[walllamp_290,floor_272]=True
    close[walllamp_290,floor_273]=True
    close[walllamp_290,ceiling_279]=True
    close[walllamp_290,bathroom_cabinet_305]=True
    close[walllamp_290,bathroom_counter_306]=True
    close[walllamp_290,sink_307]=True
    close[walllamp_290,floor_331]=True
    close[walllamp_290,floor_332]=True
    close[walllamp_290,wall_339]=True
    close[walllamp_290,wall_342]=True
    close[walllamp_290,ceiling_349]=True
    close[walllamp_290,ceiling_350]=True
    close[walllamp_290,photoframe_361]=True
    close[walllamp_290,bookshelf_372]=True
    close[walllamp_291,floor_162]=True
    close[walllamp_291,floor_163]=True
    close[walllamp_291,floor_166]=True
    close[walllamp_291,wall_169]=True
    close[walllamp_291,wall_171]=True
    close[walllamp_291,ceiling_175]=True
    close[walllamp_291,ceiling_176]=True
    close[walllamp_291,walllamp_183]=True
    close[walllamp_291,walllamp_184]=True
    close[walllamp_291,tvstand_186]=True
    close[walllamp_291,television_216]=True
    close[walllamp_291,wall_267]=True
    close[walllamp_291,wall_268]=True
    close[walllamp_291,floor_277]=True
    close[walllamp_291,floor_278]=True
    close[walllamp_291,ceiling_281]=True
    close[walllamp_291,ceiling_282]=True
    close[walllamp_291,shower_303]=True
    close[walllamp_291,curtain_304]=True
    close[curtain_293,wall_267]=True
    close[curtain_293,wall_270]=True
    close[curtain_293,floor_275]=True
    close[curtain_293,ceiling_282]=True
    close[curtain_293,ceiling_283]=True
    close[curtain_293,window_287]=True
    close[curtain_293,curtain_294]=True
    close[curtain_293,bathtub_297]=True
    close[curtain_294,wall_267]=True
    close[curtain_294,wall_270]=True
    close[curtain_294,floor_275]=True
    close[curtain_294,ceiling_282]=True
    close[curtain_294,ceiling_283]=True
    close[curtain_294,window_287]=True
    close[curtain_294,curtain_293]=True
    close[curtain_294,bathtub_297]=True
    close[bathtub_297,washing_machine_2041]=True
    close[bathtub_297,wall_266]=True
    close[bathtub_297,wall_270]=True
    close[bathtub_297,floor_274]=True
    close[bathtub_297,floor_275]=True
    close[bathtub_297,window_287]=True
    close[bathtub_297,walllamp_289]=True
    close[bathtub_297,curtain_293]=True
    close[bathtub_297,curtain_294]=True
    close[bathtub_297,wallshelf_301]=True
    close[wallshelf_301,wall_266]=True
    close[wallshelf_301,wall_270]=True
    close[wallshelf_301,ceiling_283]=True
    close[wallshelf_301,ceiling_284]=True
    close[wallshelf_301,walllamp_289]=True
    close[wallshelf_301,bathtub_297]=True
    close[toilet_302,wall_3]=True
    close[toilet_302,wall_5]=True
    close[toilet_302,floor_12]=True
    close[toilet_302,floor_13]=True
    close[toilet_302,floor_14]=True
    close[toilet_302,powersocket_48]=True
    close[toilet_302,light_49]=True
    close[toilet_302,floor_166]=True
    close[toilet_302,wall_171]=True
    close[toilet_302,walllamp_183]=True
    close[toilet_302,tvstand_186]=True
    close[toilet_302,wall_268]=True
    close[toilet_302,floor_277]=True
    close[shower_303,floor_162]=True
    close[shower_303,floor_163]=True
    close[shower_303,wall_169]=True
    close[shower_303,ceiling_175]=True
    close[shower_303,walllamp_184]=True
    close[shower_303,tvstand_186]=True
    close[shower_303,wallshelf_187]=True
    close[shower_303,wallshelf_190]=True
    close[shower_303,wallshelf_191]=True
    close[shower_303,television_216]=True
    close[shower_303,wall_267]=True
    close[shower_303,floor_278]=True
    close[shower_303,ceiling_282]=True
    close[shower_303,walllamp_291]=True
    close[shower_303,curtain_304]=True
    close[curtain_304,floor_162]=True
    close[curtain_304,floor_163]=True
    close[curtain_304,wall_169]=True
    close[curtain_304,wall_171]=True
    close[curtain_304,ceiling_175]=True
    close[curtain_304,walllamp_184]=True
    close[curtain_304,tvstand_186]=True
    close[curtain_304,television_216]=True
    close[curtain_304,wall_267]=True
    close[curtain_304,wall_268]=True
    close[curtain_304,floor_278]=True
    close[curtain_304,ceiling_282]=True
    close[curtain_304,walllamp_291]=True
    close[curtain_304,shower_303]=True
    close[bathroom_cabinet_305,wall_266]=True
    close[bathroom_cabinet_305,wall_269]=True
    close[bathroom_cabinet_305,ceiling_279]=True
    close[bathroom_cabinet_305,ceiling_284]=True
    close[bathroom_cabinet_305,walllamp_289]=True
    close[bathroom_cabinet_305,walllamp_290]=True
    close[bathroom_cabinet_305,bathroom_counter_306]=True
    close[bathroom_cabinet_305,sink_307]=True
    close[bathroom_cabinet_305,faucet_308]=True
    close[bathroom_cabinet_305,wall_339]=True
    close[bathroom_cabinet_305,photoframe_361]=True
    close[bathroom_cabinet_305,bookshelf_372]=True
    close[bathroom_counter_306,wall_266]=True
    close[bathroom_counter_306,wall_269]=True
    close[bathroom_counter_306,floor_272]=True
    close[bathroom_counter_306,floor_273]=True
    close[bathroom_counter_306,floor_274]=True
    close[bathroom_counter_306,walllamp_289]=True
    close[bathroom_counter_306,walllamp_290]=True
    close[bathroom_counter_306,bathroom_cabinet_305]=True
    close[bathroom_counter_306,sink_307]=True
    close[bathroom_counter_306,faucet_308]=True
    close[bathroom_counter_306,wall_339]=True
    close[bathroom_counter_306,photoframe_361]=True
    close[bathroom_counter_306,bookshelf_372]=True
    close[sink_307,wall_266]=True
    close[sink_307,wall_269]=True
    close[sink_307,floor_272]=True
    close[sink_307,floor_273]=True
    close[sink_307,floor_274]=True
    close[sink_307,walllamp_290]=True
    close[sink_307,bathroom_cabinet_305]=True
    close[sink_307,bathroom_counter_306]=True
    close[sink_307,faucet_308]=True
    close[faucet_308,wall_266]=True
    close[faucet_308,wall_269]=True
    close[faucet_308,floor_272]=True
    close[faucet_308,floor_273]=True
    close[faucet_308,floor_274]=True
    close[faucet_308,ceiling_279]=True
    close[faucet_308,bathroom_cabinet_305]=True
    close[faucet_308,bathroom_counter_306]=True
    close[faucet_308,sink_307]=True
    close[light_325,wall_269]=True
    close[light_325,wall_271]=True
    close[light_325,floor_272]=True
    close[light_325,floor_273]=True
    close[light_325,floor_276]=True
    close[light_325,ceiling_279]=True
    close[light_325,ceiling_280]=True
    close[light_325,doorjamb_285]=True
    close[light_325,door_286]=True
    close[light_325,floor_332]=True
    close[light_325,floor_337]=True
    close[light_325,wall_339]=True
    close[light_325,wall_345]=True
    close[light_325,ceiling_350]=True
    close[light_325,ceiling_355]=True
    close[floor_328,floor_329]=True
    close[floor_328,floor_330]=True
    close[floor_328,floor_334]=True
    close[floor_328,wall_341]=True
    close[floor_328,tablelamp_358]=True
    close[floor_328,trashcan_360]=True
    close[floor_328,bed_376]=True
    close[floor_329,floor_328]=True
    close[floor_329,floor_330]=True
    close[floor_329,floor_334]=True
    close[floor_329,wall_341]=True
    close[floor_329,tablelamp_358]=True
    close[floor_329,trashcan_360]=True
    close[floor_329,bed_376]=True
    close[floor_330,floor_328]=True
    close[floor_330,floor_329]=True
    close[floor_330,floor_331]=True
    close[floor_330,floor_333]=True
    close[floor_330,wall_340]=True
    close[floor_330,wall_341]=True
    close[floor_330,wall_342]=True
    close[floor_330,window_346]=True
    close[floor_330,tablelamp_358]=True
    close[floor_330,tablelamp_359]=True
    close[floor_330,nightstand_373]=True
    close[floor_330,bed_376]=True
    close[floor_330,curtain_390]=True
    close[floor_330,curtain_391]=True
    close[floor_330,curtain_392]=True
    close[floor_331,walllamp_290]=True
    close[floor_331,floor_330]=True
    close[floor_331,floor_332]=True
    close[floor_331,wall_342]=True
    close[floor_331,tablelamp_359]=True
    close[floor_331,bookshelf_372]=True
    close[floor_331,nightstand_373]=True
    close[floor_332,wall_269]=True
    close[floor_332,floor_272]=True
    close[floor_332,floor_273]=True
    close[floor_332,door_286]=True
    close[floor_332,walllamp_290]=True
    close[floor_332,light_325]=True
    close[floor_332,floor_331]=True
    close[floor_332,floor_333]=True
    close[floor_332,floor_337]=True
    close[floor_332,wall_339]=True
    close[floor_332,wall_342]=True
    close[floor_332,wall_345]=True
    close[floor_332,bookshelf_372]=True
    close[floor_333,floor_330]=True
    close[floor_333,floor_332]=True
    close[floor_333,floor_334]=True
    close[floor_333,floor_336]=True
    close[floor_333,bed_376]=True
    close[floor_334,floor_328]=True
    close[floor_334,floor_329]=True
    close[floor_334,floor_333]=True
    close[floor_334,floor_335]=True
    close[floor_334,wall_338]=True
    close[floor_334,wall_341]=True
    close[floor_334,wall_343]=True
    close[floor_334,trashcan_360]=True
    close[floor_334,bed_376]=True
    close[floor_334,dresser_377]=True
    close[floor_334,filing_cabinet_378]=True
    close[floor_335,wall_9]=True
    close[floor_335,floor_19]=True
    close[floor_335,door_38]=True
    close[floor_335,orchid_117]=True
    close[floor_335,tvstand_135]=True
    close[floor_335,bookshelf_137]=True
    close[floor_335,floor_334]=True
    close[floor_335,floor_336]=True
    close[floor_335,wall_343]=True
    close[floor_335,filing_cabinet_378]=True
    close[floor_335,light_384]=True
    close[floor_336,wall_10]=True
    close[floor_336,floor_18]=True
    close[floor_336,door_38]=True
    close[floor_336,orchid_117]=True
    close[floor_336,tvstand_135]=True
    close[floor_336,bookshelf_136]=True
    close[floor_336,floor_333]=True
    close[floor_336,floor_335]=True
    close[floor_336,floor_337]=True
    close[floor_336,wall_343]=True
    close[floor_336,wall_344]=True
    close[floor_336,wall_345]=True
    close[floor_336,doorjamb_356]=True
    close[floor_336,desk_375]=True
    close[floor_336,computer_379]=True
    close[floor_336,mousepad_381]=True
    close[floor_336,cpuscreen_383]=True
    close[floor_336,light_384]=True
    close[floor_337,wall_5]=True
    close[floor_337,floor_12]=True
    close[floor_337,floor_13]=True
    close[floor_337,door_38]=True
    close[floor_337,bookshelf_136]=True
    close[floor_337,wall_271]=True
    close[floor_337,floor_276]=True
    close[floor_337,doorjamb_285]=True
    close[floor_337,door_286]=True
    close[floor_337,light_325]=True
    close[floor_337,floor_332]=True
    close[floor_337,floor_336]=True
    close[floor_337,wall_345]=True
    close[floor_337,desk_375]=True
    close[floor_337,computer_379]=True
    close[floor_337,mousepad_381]=True
    close[floor_337,cpuscreen_383]=True
    close[wall_338,floor_334]=True
    close[wall_338,wall_341]=True
    close[wall_338,wall_343]=True
    close[wall_338,ceiling_352]=True
    close[wall_338,trashcan_360]=True
    close[wall_338,dresser_377]=True
    close[wall_338,filing_cabinet_378]=True
    close[wall_339,wall_269]=True
    close[wall_339,wall_271]=True
    close[wall_339,floor_272]=True
    close[wall_339,floor_273]=True
    close[wall_339,ceiling_279]=True
    close[wall_339,doorjamb_285]=True
    close[wall_339,door_286]=True
    close[wall_339,walllamp_290]=True
    close[wall_339,bathroom_cabinet_305]=True
    close[wall_339,bathroom_counter_306]=True
    close[wall_339,light_325]=True
    close[wall_339,floor_332]=True
    close[wall_339,wall_342]=True
    close[wall_339,wall_345]=True
    close[wall_339,ceiling_350]=True
    close[wall_339,photoframe_361]=True
    close[wall_339,bookshelf_372]=True
    close[wall_340,floor_330]=True
    close[wall_340,wall_341]=True
    close[wall_340,wall_342]=True
    close[wall_340,window_346]=True
    close[wall_340,ceiling_348]=True
    close[wall_340,tablelamp_358]=True
    close[wall_340,tablelamp_359]=True
    close[wall_340,nightstand_373]=True
    close[wall_340,bed_376]=True
    close[wall_340,curtain_390]=True
    close[wall_340,curtain_391]=True
    close[wall_340,curtain_392]=True
    close[wall_341,floor_328]=True
    close[wall_341,floor_329]=True
    close[wall_341,floor_330]=True
    close[wall_341,floor_334]=True
    close[wall_341,wall_338]=True
    close[wall_341,wall_340]=True
    close[wall_341,window_346]=True
    close[wall_341,ceiling_347]=True
    close[wall_341,ceiling_348]=True
    close[wall_341,ceiling_352]=True
    close[wall_341,tablelamp_358]=True
    close[wall_341,trashcan_360]=True
    close[wall_341,bed_376]=True
    close[wall_341,dresser_377]=True
    close[wall_341,curtain_390]=True
    close[wall_341,curtain_391]=True
    close[wall_342,walllamp_290]=True
    close[wall_342,floor_330]=True
    close[wall_342,floor_331]=True
    close[wall_342,floor_332]=True
    close[wall_342,wall_339]=True
    close[wall_342,wall_340]=True
    close[wall_342,window_346]=True
    close[wall_342,ceiling_348]=True
    close[wall_342,ceiling_349]=True
    close[wall_342,ceiling_350]=True
    close[wall_342,tablelamp_359]=True
    close[wall_342,photoframe_361]=True
    close[wall_342,bookshelf_372]=True
    close[wall_342,nightstand_373]=True
    close[wall_342,curtain_392]=True
    close[wall_343,wall_9]=True
    close[wall_343,wall_10]=True
    close[wall_343,floor_19]=True
    close[wall_343,ceiling_31]=True
    close[wall_343,door_38]=True
    close[wall_343,orchid_117]=True
    close[wall_343,tvstand_135]=True
    close[wall_343,bookshelf_137]=True
    close[wall_343,floor_334]=True
    close[wall_343,floor_335]=True
    close[wall_343,floor_336]=True
    close[wall_343,wall_338]=True
    close[wall_343,wall_344]=True
    close[wall_343,ceiling_352]=True
    close[wall_343,ceiling_353]=True
    close[wall_343,ceiling_354]=True
    close[wall_343,doorjamb_356]=True
    close[wall_343,dresser_377]=True
    close[wall_343,filing_cabinet_378]=True
    close[wall_343,light_384]=True
    close[wall_344,wall_5]=True
    close[wall_344,wall_9]=True
    close[wall_344,wall_10]=True
    close[wall_344,floor_18]=True
    close[wall_344,ceiling_30]=True
    close[wall_344,door_38]=True
    close[wall_344,orchid_117]=True
    close[wall_344,tvstand_135]=True
    close[wall_344,bookshelf_136]=True
    close[wall_344,floor_336]=True
    close[wall_344,wall_343]=True
    close[wall_344,wall_345]=True
    close[wall_344,ceiling_354]=True
    close[wall_344,doorjamb_356]=True
    close[wall_344,desk_375]=True
    close[wall_344,computer_379]=True
    close[wall_344,mousepad_381]=True
    close[wall_344,cpuscreen_383]=True
    close[wall_344,light_384]=True
    close[wall_345,wall_5]=True
    close[wall_345,wall_10]=True
    close[wall_345,floor_12]=True
    close[wall_345,floor_13]=True
    close[wall_345,ceiling_25]=True
    close[wall_345,door_38]=True
    close[wall_345,bookshelf_136]=True
    close[wall_345,wall_271]=True
    close[wall_345,floor_276]=True
    close[wall_345,ceiling_280]=True
    close[wall_345,doorjamb_285]=True
    close[wall_345,door_286]=True
    close[wall_345,light_325]=True
    close[wall_345,floor_332]=True
    close[wall_345,floor_336]=True
    close[wall_345,floor_337]=True
    close[wall_345,wall_339]=True
    close[wall_345,wall_344]=True
    close[wall_345,ceiling_350]=True
    close[wall_345,ceiling_354]=True
    close[wall_345,ceiling_355]=True
    close[wall_345,doorjamb_356]=True
    close[wall_345,desk_375]=True
    close[wall_345,computer_379]=True
    close[wall_345,mousepad_381]=True
    close[wall_345,cpuscreen_383]=True
    close[window_346,floor_330]=True
    close[window_346,wall_340]=True
    close[window_346,wall_341]=True
    close[window_346,wall_342]=True
    close[window_346,ceiling_348]=True
    close[window_346,tablelamp_358]=True
    close[window_346,tablelamp_359]=True
    close[window_346,nightstand_373]=True
    close[window_346,bed_376]=True
    close[window_346,curtain_390]=True
    close[window_346,curtain_391]=True
    close[window_346,curtain_392]=True
    close[ceiling_347,wall_341]=True
    close[ceiling_347,ceiling_348]=True
    close[ceiling_347,ceiling_352]=True
    close[ceiling_347,curtain_390]=True
    close[ceiling_347,curtain_391]=True
    close[ceiling_348,wall_340]=True
    close[ceiling_348,wall_341]=True
    close[ceiling_348,wall_342]=True
    close[ceiling_348,window_346]=True
    close[ceiling_348,ceiling_347]=True
    close[ceiling_348,ceiling_349]=True
    close[ceiling_348,ceiling_351]=True
    close[ceiling_348,ceilinglamp_357]=True
    close[ceiling_348,curtain_390]=True
    close[ceiling_348,curtain_391]=True
    close[ceiling_348,curtain_392]=True
    close[ceiling_349,walllamp_290]=True
    close[ceiling_349,wall_342]=True
    close[ceiling_349,ceiling_348]=True
    close[ceiling_349,ceiling_350]=True
    close[ceiling_349,photoframe_361]=True
    close[ceiling_349,bookshelf_372]=True
    close[ceiling_349,curtain_392]=True
    close[ceiling_350,wall_269]=True
    close[ceiling_350,ceiling_279]=True
    close[ceiling_350,walllamp_290]=True
    close[ceiling_350,light_325]=True
    close[ceiling_350,wall_339]=True
    close[ceiling_350,wall_342]=True
    close[ceiling_350,wall_345]=True
    close[ceiling_350,ceiling_349]=True
    close[ceiling_350,ceiling_351]=True
    close[ceiling_350,ceiling_355]=True
    close[ceiling_350,ceilinglamp_357]=True
    close[ceiling_350,photoframe_361]=True
    close[ceiling_350,bookshelf_372]=True
    close[ceiling_351,ceiling_348]=True
    close[ceiling_351,ceiling_350]=True
    close[ceiling_351,ceiling_352]=True
    close[ceiling_351,ceiling_354]=True
    close[ceiling_351,ceilinglamp_357]=True
    close[ceiling_352,wall_338]=True
    close[ceiling_352,wall_341]=True
    close[ceiling_352,wall_343]=True
    close[ceiling_352,ceiling_347]=True
    close[ceiling_352,ceiling_351]=True
    close[ceiling_352,ceiling_353]=True
    close[ceiling_352,ceilinglamp_357]=True
    close[ceiling_352,dresser_377]=True
    close[ceiling_353,wall_9]=True
    close[ceiling_353,ceiling_31]=True
    close[ceiling_353,wall_343]=True
    close[ceiling_353,ceiling_352]=True
    close[ceiling_353,ceiling_354]=True
    close[ceiling_353,light_384]=True
    close[ceiling_354,wall_10]=True
    close[ceiling_354,ceiling_30]=True
    close[ceiling_354,wall_343]=True
    close[ceiling_354,wall_344]=True
    close[ceiling_354,wall_345]=True
    close[ceiling_354,ceiling_351]=True
    close[ceiling_354,ceiling_353]=True
    close[ceiling_354,ceiling_355]=True
    close[ceiling_354,doorjamb_356]=True
    close[ceiling_354,ceilinglamp_357]=True
    close[ceiling_354,cpuscreen_383]=True
    close[ceiling_354,light_384]=True
    close[ceiling_355,wall_5]=True
    close[ceiling_355,ceiling_25]=True
    close[ceiling_355,bookshelf_136]=True
    close[ceiling_355,wall_271]=True
    close[ceiling_355,ceiling_280]=True
    close[ceiling_355,doorjamb_285]=True
    close[ceiling_355,light_325]=True
    close[ceiling_355,wall_345]=True
    close[ceiling_355,ceiling_350]=True
    close[ceiling_355,ceiling_354]=True
    close[ceiling_355,cpuscreen_383]=True
    close[doorjamb_356,wall_5]=True
    close[doorjamb_356,wall_9]=True
    close[doorjamb_356,wall_10]=True
    close[doorjamb_356,floor_18]=True
    close[doorjamb_356,ceiling_30]=True
    close[doorjamb_356,door_38]=True
    close[doorjamb_356,bookshelf_136]=True
    close[doorjamb_356,floor_336]=True
    close[doorjamb_356,wall_343]=True
    close[doorjamb_356,wall_344]=True
    close[doorjamb_356,wall_345]=True
    close[doorjamb_356,ceiling_354]=True
    close[doorjamb_356,desk_375]=True
    close[doorjamb_356,mousepad_381]=True
    close[doorjamb_356,cpuscreen_383]=True
    close[doorjamb_356,light_384]=True
    close[ceilinglamp_357,ceiling_348]=True
    close[ceilinglamp_357,ceiling_350]=True
    close[ceilinglamp_357,ceiling_351]=True
    close[ceilinglamp_357,ceiling_352]=True
    close[ceilinglamp_357,ceiling_354]=True
    close[tablelamp_358,floor_328]=True
    close[tablelamp_358,floor_329]=True
    close[tablelamp_358,floor_330]=True
    close[tablelamp_358,wall_340]=True
    close[tablelamp_358,wall_341]=True
    close[tablelamp_358,window_346]=True
    close[tablelamp_358,bed_376]=True
    close[tablelamp_358,curtain_390]=True
    close[tablelamp_358,curtain_391]=True
    close[tablelamp_359,floor_330]=True
    close[tablelamp_359,floor_331]=True
    close[tablelamp_359,wall_340]=True
    close[tablelamp_359,wall_342]=True
    close[tablelamp_359,window_346]=True
    close[tablelamp_359,nightstand_373]=True
    close[tablelamp_359,bed_376]=True
    close[tablelamp_359,curtain_390]=True
    close[tablelamp_359,curtain_391]=True
    close[tablelamp_359,curtain_392]=True
    close[trashcan_360,floor_328]=True
    close[trashcan_360,floor_329]=True
    close[trashcan_360,floor_334]=True
    close[trashcan_360,wall_338]=True
    close[trashcan_360,wall_341]=True
    close[photoframe_361,wall_269]=True
    close[photoframe_361,ceiling_279]=True
    close[photoframe_361,walllamp_290]=True
    close[photoframe_361,bathroom_cabinet_305]=True
    close[photoframe_361,bathroom_counter_306]=True
    close[photoframe_361,wall_339]=True
    close[photoframe_361,wall_342]=True
    close[photoframe_361,ceiling_349]=True
    close[photoframe_361,ceiling_350]=True
    close[photoframe_361,bookshelf_372]=True
    close[bookshelf_372,wall_269]=True
    close[bookshelf_372,floor_272]=True
    close[bookshelf_372,floor_273]=True
    close[bookshelf_372,ceiling_279]=True
    close[bookshelf_372,walllamp_290]=True
    close[bookshelf_372,bathroom_cabinet_305]=True
    close[bookshelf_372,bathroom_counter_306]=True
    close[bookshelf_372,floor_331]=True
    close[bookshelf_372,floor_332]=True
    close[bookshelf_372,wall_339]=True
    close[bookshelf_372,wall_342]=True
    close[bookshelf_372,ceiling_349]=True
    close[bookshelf_372,ceiling_350]=True
    close[bookshelf_372,photoframe_361]=True
    close[nightstand_373,floor_330]=True
    close[nightstand_373,floor_331]=True
    close[nightstand_373,wall_340]=True
    close[nightstand_373,wall_342]=True
    close[nightstand_373,window_346]=True
    close[nightstand_373,tablelamp_359]=True
    close[nightstand_373,bed_376]=True
    close[nightstand_373,curtain_390]=True
    close[nightstand_373,curtain_391]=True
    close[nightstand_373,curtain_392]=True
    close[desk_375,wall_5]=True
    close[desk_375,wall_10]=True
    close[desk_375,floor_12]=True
    close[desk_375,floor_13]=True
    close[desk_375,floor_18]=True
    close[desk_375,door_38]=True
    close[desk_375,bookshelf_136]=True
    close[desk_375,wall_271]=True
    close[desk_375,doorjamb_285]=True
    close[desk_375,door_286]=True
    close[desk_375,floor_336]=True
    close[desk_375,floor_337]=True
    close[desk_375,wall_344]=True
    close[desk_375,wall_345]=True
    close[desk_375,doorjamb_356]=True
    close[desk_375,computer_379]=True
    close[desk_375,mousepad_381]=True
    close[desk_375,cpuscreen_383]=True
    close[desk_375,light_384]=True
    close[bed_376,floor_328]=True
    close[bed_376,floor_329]=True
    close[bed_376,floor_330]=True
    close[bed_376,floor_333]=True
    close[bed_376,floor_334]=True
    close[bed_376,wall_340]=True
    close[bed_376,wall_341]=True
    close[bed_376,window_346]=True
    close[bed_376,tablelamp_358]=True
    close[bed_376,tablelamp_359]=True
    close[bed_376,nightstand_373]=True
    close[bed_376,curtain_390]=True
    close[bed_376,curtain_391]=True
    close[bed_376,curtain_392]=True
    close[dresser_377,floor_334]=True
    close[dresser_377,wall_338]=True
    close[dresser_377,wall_341]=True
    close[dresser_377,wall_343]=True
    close[dresser_377,ceiling_352]=True
    close[dresser_377,filing_cabinet_378]=True
    close[filing_cabinet_378,wall_9]=True
    close[filing_cabinet_378,wall_11]=True
    close[filing_cabinet_378,bookshelf_137]=True
    close[filing_cabinet_378,floor_334]=True
    close[filing_cabinet_378,floor_335]=True
    close[filing_cabinet_378,wall_338]=True
    close[filing_cabinet_378,wall_343]=True
    close[filing_cabinet_378,dresser_377]=True
    close[computer_379,wall_5]=True
    close[computer_379,wall_10]=True
    close[computer_379,floor_12]=True
    close[computer_379,floor_13]=True
    close[computer_379,floor_18]=True
    close[computer_379,bookshelf_136]=True
    close[computer_379,doorjamb_285]=True
    close[computer_379,door_286]=True
    close[computer_379,floor_336]=True
    close[computer_379,floor_337]=True
    close[computer_379,wall_344]=True
    close[computer_379,wall_345]=True
    close[computer_379,desk_375]=True
    close[computer_379,mousepad_381]=True
    close[computer_379,cpuscreen_383]=True
    close[mousepad_381,wall_5]=True
    close[mousepad_381,wall_10]=True
    close[mousepad_381,floor_12]=True
    close[mousepad_381,floor_13]=True
    close[mousepad_381,floor_18]=True
    close[mousepad_381,door_38]=True
    close[mousepad_381,bookshelf_136]=True
    close[mousepad_381,floor_336]=True
    close[mousepad_381,floor_337]=True
    close[mousepad_381,wall_344]=True
    close[mousepad_381,wall_345]=True
    close[mousepad_381,doorjamb_356]=True
    close[mousepad_381,desk_375]=True
    close[mousepad_381,computer_379]=True
    close[mousepad_381,cpuscreen_383]=True
    close[mousepad_381,light_384]=True
    close[cpuscreen_383,wall_5]=True
    close[cpuscreen_383,wall_10]=True
    close[cpuscreen_383,floor_12]=True
    close[cpuscreen_383,floor_13]=True
    close[cpuscreen_383,floor_18]=True
    close[cpuscreen_383,ceiling_25]=True
    close[cpuscreen_383,ceiling_30]=True
    close[cpuscreen_383,door_38]=True
    close[cpuscreen_383,bookshelf_136]=True
    close[cpuscreen_383,floor_336]=True
    close[cpuscreen_383,floor_337]=True
    close[cpuscreen_383,wall_344]=True
    close[cpuscreen_383,wall_345]=True
    close[cpuscreen_383,ceiling_354]=True
    close[cpuscreen_383,ceiling_355]=True
    close[cpuscreen_383,doorjamb_356]=True
    close[cpuscreen_383,desk_375]=True
    close[cpuscreen_383,computer_379]=True
    close[cpuscreen_383,mousepad_381]=True
    close[light_384,wall_9]=True
    close[light_384,wall_10]=True
    close[light_384,floor_18]=True
    close[light_384,floor_19]=True
    close[light_384,ceiling_30]=True
    close[light_384,ceiling_31]=True
    close[light_384,door_38]=True
    close[light_384,orchid_117]=True
    close[light_384,tvstand_135]=True
    close[light_384,floor_335]=True
    close[light_384,floor_336]=True
    close[light_384,wall_343]=True
    close[light_384,wall_344]=True
    close[light_384,ceiling_353]=True
    close[light_384,ceiling_354]=True
    close[light_384,doorjamb_356]=True
    close[light_384,desk_375]=True
    close[light_384,mousepad_381]=True
    close[curtain_390,floor_330]=True
    close[curtain_390,wall_340]=True
    close[curtain_390,wall_341]=True
    close[curtain_390,window_346]=True
    close[curtain_390,ceiling_347]=True
    close[curtain_390,ceiling_348]=True
    close[curtain_390,tablelamp_358]=True
    close[curtain_390,tablelamp_359]=True
    close[curtain_390,nightstand_373]=True
    close[curtain_390,bed_376]=True
    close[curtain_390,curtain_391]=True
    close[curtain_390,curtain_392]=True
    close[curtain_391,floor_330]=True
    close[curtain_391,wall_340]=True
    close[curtain_391,wall_341]=True
    close[curtain_391,window_346]=True
    close[curtain_391,ceiling_347]=True
    close[curtain_391,ceiling_348]=True
    close[curtain_391,tablelamp_358]=True
    close[curtain_391,tablelamp_359]=True
    close[curtain_391,nightstand_373]=True
    close[curtain_391,bed_376]=True
    close[curtain_391,curtain_390]=True
    close[curtain_391,curtain_392]=True
    close[curtain_392,floor_330]=True
    close[curtain_392,wall_340]=True
    close[curtain_392,wall_342]=True
    close[curtain_392,window_346]=True
    close[curtain_392,ceiling_348]=True
    close[curtain_392,ceiling_349]=True
    close[curtain_392,tablelamp_359]=True
    close[curtain_392,nightstand_373]=True
    close[curtain_392,bed_376]=True
    close[curtain_392,curtain_390]=True
    close[curtain_392,curtain_391]=True
    close[food_orange_2008,kitchen_counter_128]=True
    facing[wall_3,television_216]=True
    facing[wall_6,television_216]=True
    facing[doorjamb_37,television_216]=True
    facing[floor_162,television_216]=True
    facing[floor_163,television_216]=True
    facing[floor_168,television_216]=True
    facing[wall_169,television_216]=True
    facing[wall_171,television_216]=True
    facing[wall_173,television_216]=True
    facing[ceiling_175,television_216]=True
    facing[ceiling_176,television_216]=True
    facing[ceiling_177,television_216]=True
    facing[ceiling_178,television_216]=True
    facing[window_181,television_216]=True
    facing[ceilinglamp_185,television_216]=True
    facing[wallshelf_187,television_216]=True
    facing[bookshelf_189,television_216]=True
    facing[wallshelf_190,television_216]=True
    facing[wallshelf_191,television_216]=True
    facing[curtain_197,television_216]=True
    facing[curtain_198,television_216]=True
    facing[curtain_199,television_216]=True
    facing[orchid_200,television_216]=True
    facing[photoframe_210,television_216]=True
    facing[light_217,television_216]=True
    facing[powersocket_218,television_216]=True
    facing[floor_272,computer_379]=True
    facing[floor_273,computer_379]=True
    facing[floor_332,computer_379]=True
    facing[floor_333,computer_379]=True
    facing[floor_336,computer_379]=True
    facing[floor_337,computer_379]=True
    facing[wall_339,computer_379]=True
    facing[wall_345,computer_379]=True
    facing[ceiling_350,computer_379]=True
    facing[ceiling_351,computer_379]=True
    facing[ceiling_354,computer_379]=True
    facing[bookshelf_372,computer_379]=True
    #relations_end

    #exploration
    unknown[keyboard_2111]=True
    unknown[mouse_2112]=True
    unknown[clothes_pants_2113]=True
    unknown[clothes_shirt_2114]=True
    unknown[clothes_socks_2115]=True
    unknown[clothes_skirt_2116]=True
    unknown[iron_2117]=True
    unknown[chair_2118]=True
    unknown[basket_for_clothes_2040]=True
    unknown[food_steak_2042]=True
    unknown[food_apple_2043]=True
    unknown[food_bacon_2044]=True
    unknown[food_banana_2045]=True
    unknown[food_cake_2046]=True
    unknown[food_carrot_2047]=True
    unknown[food_cereal_2048]=True
    unknown[food_cheese_2049]=True
    unknown[food_chicken_2050]=True
    unknown[food_dessert_2051]=True
    unknown[food_donut_2052]=True
    unknown[food_egg_2053]=True
    unknown[food_fish_2054]=True
    unknown[food_food_2055]=True
    unknown[food_fruit_2056]=True
    unknown[food_hamburger_2057]=True
    unknown[food_ice_cream_2058]=True
    unknown[food_jam_2059]=True
    unknown[food_kiwi_2060]=True
    unknown[food_lemon_2061]=True
    unknown[food_noodles_2062]=True
    unknown[food_oatmeal_2063]=True
    unknown[food_peanut_butter_2064]=True
    unknown[food_pizza_2065]=True
    unknown[food_potato_2066]=True
    unknown[food_rice_2067]=True
    unknown[food_salt_2068]=True
    unknown[food_snack_2069]=True
    unknown[food_sugar_2070]=True
    unknown[food_turkey_2071]=True
    unknown[food_vegetable_2072]=True
    unknown[dry_pasta_2073]=True
    unknown[milk_2074]=True
    unknown[clothes_dress_2075]=True
    unknown[clothes_hat_2076]=True
    unknown[clothes_gloves_2077]=True
    unknown[clothes_jacket_2078]=True
    unknown[clothes_scarf_2079]=True
    unknown[remote_control_2081]=True
    unknown[cat_2082]=True
    unknown[towel_2083]=True
    unknown[cd_player_2084]=True
    unknown[dvd_player_2085]=True
    unknown[headset_2086]=True
    unknown[cup_2087]=True
    unknown[cup_2088]=True
    unknown[cup_2089]=True
    unknown[book_2091]=True
    unknown[book_2092]=True
    unknown[pot_2093]=True
    unknown[vacuum_cleaner_2094]=True
    unknown[bowl_2095]=True
    unknown[bowl_2096]=True
    unknown[bowl_2097]=True
    unknown[cleaning_solution_2098]=True
    unknown[cd_2100]=True
    unknown[sauce_2101]=True
    unknown[oil_2102]=True
    unknown[fork_2103]=True
    unknown[fork_2104]=True
    unknown[plate_2105]=True
    unknown[fryingpan_2107]=True
    unknown[detergent_2108]=True
    unknown[phone_47]=True
    unknown[pot_54]=True
    unknown[mat_114]=True
    unknown[mat_115]=True
    unknown[drawing_118]=True
    unknown[chair_138]=True
    unknown[tray_142]=True
    unknown[pillow_195]=True
    unknown[drawing_196]=True
    unknown[mat_201]=True
    unknown[mat_237]=True
    unknown[drawing_238]=True
    unknown[pillow_239]=True
    unknown[pillow_240]=True
    unknown[chair_263]=True
    unknown[mat_292]=True
    unknown[drawing_296]=True
    unknown[towel_rack_298]=True
    unknown[towel_rack_299]=True
    unknown[towel_rack_300]=True
    unknown[pillow_368]=True
    unknown[pillow_370]=True
    unknown[chair_374]=True
    unknown[mouse_380]=True
    unknown[keyboard_382]=True
    unknown[mat_386]=True
    unknown[drawing_387]=True
    unknown[drawing_388]=True
    unknown[drawing_389]=True
    unknown[dvd_player_2000]=True
    unknown[shoes_2001]=True
    unknown[alcohol_2002]=True
    unknown[mouse_2003]=True
    unknown[coin_2004]=True
    unknown[oil_2005]=True
    unknown[cup_2006]=True
    unknown[stereo_2007]=True
    unknown[bills_2009]=True
    unknown[novel_2010]=True
    unknown[homework_2011]=True
    unknown[needle_2012]=True
    unknown[glue_2013]=True
    unknown[napkin_2014]=True
    unknown[laptop_2015]=True
    unknown[food_bread_2016]=True
    unknown[tea_bag_2017]=True
    unknown[food_butter_2018]=True
    unknown[video_game_controller_2019]=True
    unknown[crayon_2020]=True
    unknown[dough_2021]=True
    unknown[clothes_underwear_2022]=True
    unknown[box_2023]=True
    unknown[needle_2024]=True
    unknown[laser_pointer_2025]=True
    unknown[food_onion_2026]=True
    unknown[console_2027]=True
    unknown[tape_2028]=True
    unknown[after_shave_2029]=True
    unknown[crayon_2030]=True
    unknown[stamp_2031]=True
    unknown[blender_2032]=True
    unknown[check_2033]=True
    unknown[juice_2034]=True
    unknown[coffee_filter_2035]=True
    unknown[knife_2036]=True
    unknown[soap_2037]=True
    unknown[soap_2038]=True
    unknown[pajamas_2039]=True
    #exploration_end

    #id
    id[keyboard_2111]=2111
    id[mouse_2112]=2112
    id[clothes_pants_2113]=2113
    id[clothes_shirt_2114]=2114
    id[clothes_socks_2115]=2115
    id[clothes_skirt_2116]=2116
    id[iron_2117]=2117
    id[chair_2118]=2118
    id[basket_for_clothes_2040]=2040
    id[washing_machine_2041]=2041
    id[food_steak_2042]=2042
    id[food_apple_2043]=2043
    id[food_bacon_2044]=2044
    id[food_banana_2045]=2045
    id[food_cake_2046]=2046
    id[food_carrot_2047]=2047
    id[food_cereal_2048]=2048
    id[food_cheese_2049]=2049
    id[food_chicken_2050]=2050
    id[food_dessert_2051]=2051
    id[food_donut_2052]=2052
    id[food_egg_2053]=2053
    id[food_fish_2054]=2054
    id[food_food_2055]=2055
    id[food_fruit_2056]=2056
    id[food_hamburger_2057]=2057
    id[food_ice_cream_2058]=2058
    id[food_jam_2059]=2059
    id[food_kiwi_2060]=2060
    id[food_lemon_2061]=2061
    id[food_noodles_2062]=2062
    id[food_oatmeal_2063]=2063
    id[food_peanut_butter_2064]=2064
    id[food_pizza_2065]=2065
    id[food_potato_2066]=2066
    id[food_rice_2067]=2067
    id[food_salt_2068]=2068
    id[food_snack_2069]=2069
    id[food_sugar_2070]=2070
    id[food_turkey_2071]=2071
    id[food_vegetable_2072]=2072
    id[dry_pasta_2073]=2073
    id[milk_2074]=2074
    id[clothes_dress_2075]=2075
    id[clothes_hat_2076]=2076
    id[clothes_gloves_2077]=2077
    id[clothes_jacket_2078]=2078
    id[clothes_scarf_2079]=2079
    id[cutting_board_2080]=2080
    id[remote_control_2081]=2081
    id[cat_2082]=2082
    id[towel_2083]=2083
    id[cd_player_2084]=2084
    id[dvd_player_2085]=2085
    id[headset_2086]=2086
    id[cup_2087]=2087
    id[cup_2088]=2088
    id[cup_2089]=2089
    id[stove_2090]=2090
    id[book_2091]=2091
    id[book_2092]=2092
    id[pot_2093]=2093
    id[vacuum_cleaner_2094]=2094
    id[bowl_2095]=2095
    id[bowl_2096]=2096
    id[bowl_2097]=2097
    id[cleaning_solution_2098]=2098
    id[ironing_board_2099]=2099
    id[cd_2100]=2100
    id[sauce_2101]=2101
    id[oil_2102]=2102
    id[fork_2103]=2103
    id[fork_2104]=2104
    id[plate_2105]=2105
    id[spectacles_2106]=2106
    id[fryingpan_2107]=2107
    id[detergent_2108]=2108
    id[window_2109]=2109
    id[computer_2110]=2110
    id[dining_room_1]=1
    id[wall_2]=2
    id[wall_3]=3
    id[wall_4]=4
    id[wall_5]=5
    id[wall_6]=6
    id[wall_7]=7
    id[wall_8]=8
    id[wall_9]=9
    id[wall_10]=10
    id[wall_11]=11
    id[floor_12]=12
    id[floor_13]=13
    id[floor_14]=14
    id[floor_15]=15
    id[floor_16]=16
    id[floor_17]=17
    id[floor_18]=18
    id[floor_19]=19
    id[floor_20]=20
    id[floor_21]=21
    id[floor_22]=22
    id[floor_23]=23
    id[floor_24]=24
    id[ceiling_25]=25
    id[ceiling_26]=26
    id[ceiling_27]=27
    id[ceiling_28]=28
    id[ceiling_29]=29
    id[ceiling_30]=30
    id[ceiling_31]=31
    id[ceiling_32]=32
    id[ceiling_33]=33
    id[ceiling_34]=34
    id[ceiling_35]=35
    id[ceiling_36]=36
    id[doorjamb_37]=37
    id[door_38]=38
    id[doorjamb_39]=39
    id[window_40]=40
    id[ceilinglamp_41]=41
    id[ceilinglamp_42]=42
    id[ceilinglamp_43]=43
    id[walllamp_44]=44
    id[walllamp_45]=45
    id[walllamp_46]=46
    id[phone_47]=47
    id[powersocket_48]=48
    id[light_49]=49
    id[knifeblock_52]=52
    id[pot_54]=54
    id[photoframe_102]=102
    id[mat_114]=114
    id[mat_115]=115
    id[orchid_117]=117
    id[drawing_118]=118
    id[curtain_119]=119
    id[curtain_120]=120
    id[curtain_121]=121
    id[bench_122]=122
    id[table_123]=123
    id[bench_124]=124
    id[bench_125]=125
    id[bench_126]=126
    id[table_127]=127
    id[kitchen_counter_128]=128
    id[kitchen_counter_129]=129
    id[cupboard_130]=130
    id[cupboard_131]=131
    id[kitchen_counter_132]=132
    id[sink_133]=133
    id[faucet_134]=134
    id[tvstand_135]=135
    id[bookshelf_136]=136
    id[bookshelf_137]=137
    id[chair_138]=138
    id[stovefan_139]=139
    id[fridge_140]=140
    id[oven_141]=141
    id[tray_142]=142
    id[dishwasher_143]=143
    id[toaster_144]=144
    id[coffe_maker_147]=147
    id[microwave_149]=149
    id[home_office_161]=161
    id[floor_162]=162
    id[floor_163]=163
    id[floor_164]=164
    id[floor_165]=165
    id[floor_166]=166
    id[floor_167]=167
    id[floor_168]=168
    id[wall_169]=169
    id[wall_170]=170
    id[wall_171]=171
    id[wall_172]=172
    id[wall_173]=173
    id[wall_174]=174
    id[ceiling_175]=175
    id[ceiling_176]=176
    id[ceiling_177]=177
    id[ceiling_178]=178
    id[ceiling_179]=179
    id[ceiling_180]=180
    id[window_181]=181
    id[doorjamb_182]=182
    id[walllamp_183]=183
    id[walllamp_184]=184
    id[ceilinglamp_185]=185
    id[tvstand_186]=186
    id[wallshelf_187]=187
    id[bookshelf_188]=188
    id[bookshelf_189]=189
    id[wallshelf_190]=190
    id[wallshelf_191]=191
    id[couch_192]=192
    id[table_193]=193
    id[pillow_195]=195
    id[drawing_196]=196
    id[curtain_197]=197
    id[curtain_198]=198
    id[curtain_199]=199
    id[orchid_200]=200
    id[mat_201]=201
    id[photoframe_210]=210
    id[television_216]=216
    id[light_217]=217
    id[powersocket_218]=218
    id[bedroom_220]=220
    id[floor_221]=221
    id[floor_222]=222
    id[floor_223]=223
    id[floor_224]=224
    id[floor_225]=225
    id[ceiling_226]=226
    id[ceiling_227]=227
    id[ceiling_228]=228
    id[ceiling_229]=229
    id[wall_230]=230
    id[wall_231]=231
    id[wall_232]=232
    id[wall_233]=233
    id[door_234]=234
    id[ceilinglamp_235]=235
    id[tablelamp_236]=236
    id[mat_237]=237
    id[drawing_238]=238
    id[pillow_239]=239
    id[pillow_240]=240
    id[photoframe_246]=246
    id[light_258]=258
    id[powersocket_259]=259
    id[bookshelf_260]=260
    id[desk_261]=261
    id[nightstand_262]=262
    id[chair_263]=263
    id[bed_264]=264
    id[bathroom_265]=265
    id[wall_266]=266
    id[wall_267]=267
    id[wall_268]=268
    id[wall_269]=269
    id[wall_270]=270
    id[wall_271]=271
    id[floor_272]=272
    id[floor_273]=273
    id[floor_274]=274
    id[floor_275]=275
    id[floor_276]=276
    id[floor_277]=277
    id[floor_278]=278
    id[ceiling_279]=279
    id[ceiling_280]=280
    id[ceiling_281]=281
    id[ceiling_282]=282
    id[ceiling_283]=283
    id[ceiling_284]=284
    id[doorjamb_285]=285
    id[door_286]=286
    id[window_287]=287
    id[ceilinglamp_288]=288
    id[walllamp_289]=289
    id[walllamp_290]=290
    id[walllamp_291]=291
    id[mat_292]=292
    id[curtain_293]=293
    id[curtain_294]=294
    id[drawing_296]=296
    id[bathtub_297]=297
    id[towel_rack_298]=298
    id[towel_rack_299]=299
    id[towel_rack_300]=300
    id[wallshelf_301]=301
    id[toilet_302]=302
    id[shower_303]=303
    id[curtain_304]=304
    id[bathroom_cabinet_305]=305
    id[bathroom_counter_306]=306
    id[sink_307]=307
    id[faucet_308]=308
    id[light_325]=325
    id[bedroom_327]=327
    id[floor_328]=328
    id[floor_329]=329
    id[floor_330]=330
    id[floor_331]=331
    id[floor_332]=332
    id[floor_333]=333
    id[floor_334]=334
    id[floor_335]=335
    id[floor_336]=336
    id[floor_337]=337
    id[wall_338]=338
    id[wall_339]=339
    id[wall_340]=340
    id[wall_341]=341
    id[wall_342]=342
    id[wall_343]=343
    id[wall_344]=344
    id[wall_345]=345
    id[window_346]=346
    id[ceiling_347]=347
    id[ceiling_348]=348
    id[ceiling_349]=349
    id[ceiling_350]=350
    id[ceiling_351]=351
    id[ceiling_352]=352
    id[ceiling_353]=353
    id[ceiling_354]=354
    id[ceiling_355]=355
    id[doorjamb_356]=356
    id[ceilinglamp_357]=357
    id[tablelamp_358]=358
    id[tablelamp_359]=359
    id[trashcan_360]=360
    id[photoframe_361]=361
    id[pillow_368]=368
    id[pillow_370]=370
    id[bookshelf_372]=372
    id[nightstand_373]=373
    id[chair_374]=374
    id[desk_375]=375
    id[bed_376]=376
    id[dresser_377]=377
    id[filing_cabinet_378]=378
    id[computer_379]=379
    id[mouse_380]=380
    id[mousepad_381]=381
    id[keyboard_382]=382
    id[cpuscreen_383]=383
    id[light_384]=384
    id[mat_386]=386
    id[drawing_387]=387
    id[drawing_388]=388
    id[drawing_389]=389
    id[curtain_390]=390
    id[curtain_391]=391
    id[curtain_392]=392
    id[dvd_player_2000]=2000
    id[shoes_2001]=2001
    id[alcohol_2002]=2002
    id[mouse_2003]=2003
    id[coin_2004]=2004
    id[oil_2005]=2005
    id[cup_2006]=2006
    id[stereo_2007]=2007
    id[food_orange_2008]=2008
    id[bills_2009]=2009
    id[novel_2010]=2010
    id[homework_2011]=2011
    id[needle_2012]=2012
    id[glue_2013]=2013
    id[napkin_2014]=2014
    id[laptop_2015]=2015
    id[food_bread_2016]=2016
    id[tea_bag_2017]=2017
    id[food_butter_2018]=2018
    id[video_game_controller_2019]=2019
    id[crayon_2020]=2020
    id[dough_2021]=2021
    id[clothes_underwear_2022]=2022
    id[box_2023]=2023
    id[needle_2024]=2024
    id[laser_pointer_2025]=2025
    id[food_onion_2026]=2026
    id[console_2027]=2027
    id[tape_2028]=2028
    id[after_shave_2029]=2029
    id[crayon_2030]=2030
    id[stamp_2031]=2031
    id[blender_2032]=2032
    id[check_2033]=2033
    id[juice_2034]=2034
    id[coffee_filter_2035]=2035
    id[knife_2036]=2036
    id[soap_2037]=2037
    id[soap_2038]=2038
    id[pajamas_2039]=2039
    #id_end

    #size
    #size_end

#exp_behavior

behavior find_pot_54_around_cupboard_131(pot:item):
    goal: not unknown(pot)
    body:
        assert is_pot(pot)
        bind cupboard_instance:item where:
            is_cupboard(cupboard_instance) and id[cupboard_instance]==131
        achieve close_char(char,cupboard_instance)
        if can_open(cupboard_instance):
            achieve_once open(cupboard_instance)
            exp(pot,cupboard_instance)
        else:
            exp(pot,cupboard_instance)
    eff:
        unknown[pot]=False
        close[pot,cupboard_instance]=True
        close[cupboard_instance,pot]=True
    

behavior find_fryingpan_2107_around_cupboard_131(fryingpan:item):
    goal: not unknown(fryingpan)
    body:
        assert is_fryingpan(fryingpan)
        bind cupboard_instance:item where:
            is_cupboard(cupboard_instance) and id[cupboard_instance]==131
        achieve close_char(char,cupboard_instance)
        if can_open(cupboard_instance):
            achieve_once open(cupboard_instance)
            exp(fryingpan,cupboard_instance)
        else:
            exp(fryingpan,cupboard_instance)
    eff:
        unknown[fryingpan]=False
        close[fryingpan,cupboard_instance]=True
        close[cupboard_instance,fryingpan]=True
    

behavior find_food_turkey_2071_around_fridge_140(food_turkey:item):
    goal: not unknown(food_turkey)
    body:
        assert is_food_turkey(food_turkey)
        bind fridge_instance:item where:
            is_fridge(fridge_instance) and id[fridge_instance]==140
        achieve close_char(char,fridge_instance)
        if can_open(fridge_instance):
            achieve_once open(fridge_instance)
            exp(food_turkey,fridge_instance)
        else:
            exp(food_turkey,fridge_instance)
    eff:
        unknown[food_turkey]=False
        close[food_turkey,fridge_instance]=True
        close[fridge_instance,food_turkey]=True
    

behavior find_dry_pasta_2073_around_cupboard_131(dry_pasta:item):
    goal: not unknown(dry_pasta)
    body:
        assert is_dry_pasta(dry_pasta)
        bind cupboard_instance:item where:
            is_cupboard(cupboard_instance) and id[cupboard_instance]==131
        achieve close_char(char,cupboard_instance)
        if can_open(cupboard_instance):
            achieve_once open(cupboard_instance)
            exp(dry_pasta,cupboard_instance)
        else:
            exp(dry_pasta,cupboard_instance)
    eff:
        unknown[dry_pasta]=False
        close[dry_pasta,cupboard_instance]=True
        close[cupboard_instance,dry_pasta]=True
    

#exp_behavior_end

#goal_representation
 
def has_faucet(sink:item):
    # Determine whether the sink has a faucet
    symbol has_faucet=exists faucet:item: is_faucet(faucet) and close(faucet,sink)
    return has_faucet

behavior boil_pasta(pasta:item, pot:item, stove:item):
    body:
        achieve inside(pasta, pot)
        achieve on(pot, stove)
        achieve is_on(stove)
        # Boil the pasta by placing it in the pot and heating it on the stove

behavior cook_chicken(chicken:item, fryingpan:item, stove:item):
    body:
        achieve inside(chicken, fryingpan)
        achieve on(fryingpan, stove)
        achieve is_on(stove)
        # Cook the chicken by placing it in the frying pan and heating it on the stove

behavior __goal__():
    body:
        bind pot: item where:
            is_pot(pot)
        # Select a pot for boiling pasta

        bind fryingpan: item where:
            is_fryingpan(fryingpan)
        # Select a frying pan for cooking chicken

        bind stove: item where:
            is_stove(stove)
        # Select a stove for both boiling pasta and cooking chicken

        bind pasta: item where:
            is_dry_pasta(pasta)
        # Select the dry pasta

        bind chicken: item where:
            is_food_chicken(chicken)
        # Select the chicken

        boil_pasta(pasta, pot, stove)
        cook_chicken(chicken, fryingpan, stove)

#goal_representation_end
