problem "agent-problem"
domain "virtualhome_partial.cdl"

objects:
  A, B, C, D: Object

init:
  is_object[A] = True
  is_object[B] = True
  is_container[C] = True
  is_container[D] = True

  can_contain[C, A] = True
  can_contain[D, A] = True
  can_contain[C, B] = True # B can only be contained in C but not D

behavior __goal__():
  body:
    achieve contained_in_something(A)
    achieve contained_in_something(B)