problem "kitchen-problem"
domain "kitchen.cdl"

#!pragma planner_is_goal_serializable=False
#!pragma planner_is_goal_ordered=True
#!pragma planner_always_commit_skeleton=True

objects:
  tomato_1:item
  tomato_2:item
  tomato_3:item
  tomato_4:item
  egg_5:item
  egg_6:item
  egg_7:item
  egg_8:item
  oil_9:item
  sugar_10:item
  pan_11:item
  salt_12:item
  bowl_13:item
  bowl_14:item
  bowl_15:item
  bowl_16:item
  knife_17:item
  fridge_18:item
  stove_19:item
  sink_20:item
  faucet_21:item
  spatula_22:item
  countertop_23:item
  water_24:item
  pepper_25:item

init:
    is_tomato[tomato_1]=True
    is_tomato[tomato_2]=True
    is_tomato[tomato_3]=True
    is_tomato[tomato_4]=True
    is_egg[egg_5]=True
    is_egg[egg_6]=True
    is_egg[egg_7]=True
    is_egg[egg_8]=True
    is_oil[oil_9]=True
    is_sugar[sugar_10]=True
    is_pan[pan_11]=True
    is_salt[salt_12]=True
    is_bowl[bowl_13]=True
    is_bowl[bowl_14]=True
    is_bowl[bowl_15]=True
    is_bowl[bowl_16]=True
    is_knife[knife_17]=True
    is_fridge[fridge_18]=True
    is_stove[stove_19]=True
    is_sink[sink_20]=True
    is_faucet[faucet_21]=True
    is_spatula[spatula_22]=True
    is_countertop[countertop_23]=True
    is_water[water_24]=True
    is_pepper[pepper_25]=True


    is_off[stove_19]=True
    is_on[stove_19]=False
    is_off[faucet_21]=True
    is_on[faucet_21]=False
    open[fridge_18]=False
    closed[fridge_18]=True
    dirty[pan_11]=False
    clean[pan_11]=True
    dirty[bowl_13]=False
    clean[bowl_13]=True
    dirty[bowl_14]=False
    clean[bowl_14]=True
    dirty[bowl_15]=False
    clean[bowl_15]=True
    dirty[bowl_16]=False
    clean[bowl_16]=True
    dirty[tomato_1]=True
    clean[tomato_1]=False
    dirty[tomato_2]=True
    clean[tomato_2]=False
    dirty[tomato_3]=True
    clean[tomato_3]=False
    dirty[tomato_4]=True
    clean[tomato_4]=False
    sliced[tomato_1]=False
    sliced[tomato_2]=False
    sliced[tomato_3]=False
    sliced[tomato_4]=False
    peeled[egg_5]=False
    peeled[egg_6]=False
    peeled[egg_7]=False
    peeled[egg_8]=False
    peeled[tomato_1]=False
    peeled[tomato_2]=False
    peeled[tomato_3]=False
    peeled[tomato_4]=False
    raw[egg_5]=True
    cooked[egg_5]=False
    raw[egg_6]=True
    cooked[egg_6]=False
    raw[egg_7]=True
    cooked[egg_7]=False
    raw[egg_8]=True
    cooked[egg_8]=False
    raw[tomato_1]=True
    cooked[tomato_1]=False
    raw[tomato_2]=True
    cooked[tomato_2]=False
    raw[tomato_3]=True
    cooked[tomato_3]=False
    raw[tomato_4]=True
    cooked[tomato_4]=False
    heated[pan_11]=False
    mixed[pan_11]=False

    surfaces[countertop_23]=True
    surfaces[stove_19]=True
    grabbable[tomato_1]=True
    grabbable[tomato_2]=True
    grabbable[tomato_3]=True
    grabbable[tomato_4]=True
    grabbable[egg_5]=True
    grabbable[egg_6]=True
    grabbable[egg_7]=True
    grabbable[egg_8]=True
    grabbable[oil_9]=True
    grabbable[sugar_10]=True
    grabbable[pan_11]=True
    grabbable[salt_12]=True
    grabbable[bowl_13]=True
    grabbable[bowl_14]=True
    grabbable[bowl_15]=True
    grabbable[bowl_16]=True
    grabbable[knife_17]=True
    grabbable[spatula_22]=True
    recipient[bowl_13]=True
    recipient[bowl_14]=True
    recipient[bowl_15]=True
    recipient[bowl_16]=True
    recipient[pan_11]=True
    recipient[sink_20]=True
    recipient[fridge_18]=True
    cuttable[tomato_1]=True
    cuttable[tomato_2]=True
    cuttable[tomato_3]=True
    cuttable[tomato_4]=True
    containers[fridge_18]=True
    containers[bowl_13]=True
    containers[bowl_14]=True
    containers[bowl_15]=True
    containers[bowl_16]=True
    containers[pan_11]=True
    containers[sink_20]=True
    peelable[tomato_1]=True
    peelable[tomato_2]=True
    peelable[tomato_3]=True
    peelable[tomato_4]=True
    can_open[fridge_18]=True
    has_switch[stove_19]=True
    has_switch[faucet_21]=True
    storable[countertop_23]=True

    inside[tomato_1,fridge_18]=True
    inside[tomato_2,fridge_18]=True
    inside[tomato_3,fridge_18]=True
    inside[tomato_4,fridge_18]=True
    close[tomato_1,fridge_18]=True
    close[tomato_2,fridge_18]=True
    close[tomato_3,fridge_18]=True
    close[tomato_4,fridge_18]=True
    close[fridge_18,tomato_1]=True
    close[fridge_18,tomato_2]=True
    close[fridge_18,tomato_3]=True
    close[fridge_18,tomato_4]=True
    inside[egg_5,fridge_18]=True
    inside[egg_6,fridge_18]=True
    inside[egg_7,fridge_18]=True
    inside[egg_8,fridge_18]=True
    close[egg_5,fridge_18]=True
    close[egg_6,fridge_18]=True
    close[egg_7,fridge_18]=True
    close[egg_8,fridge_18]=True
    close[fridge_18,egg_5]=True
    close[fridge_18,egg_6]=True
    close[fridge_18,egg_7]=True
    close[fridge_18,egg_8]=True

    on[pan_11,countertop_23]=True
    close[pan_11,countertop_23]=True
    close[countertop_23,pan_11]=True

    on[faucet_21,sink_20]=True
    close[faucet_21,sink_20]=True
    close[sink_20,faucet_21]=True
    on[bowl_13,countertop_23]=True
    close[bowl_13,countertop_23]=True
    close[countertop_23,bowl_13]=True
    on[bowl_14,countertop_23]=True
    close[bowl_14,countertop_23]=True
    close[countertop_23,bowl_14]=True
    on[bowl_15,countertop_23]=True
    close[bowl_15,countertop_23]=True
    close[countertop_23,bowl_15]=True
    on[bowl_16,countertop_23]=True
    close[bowl_16,countertop_23]=True
    close[countertop_23,bowl_16]=True
    inside[spatula_22,pan_11]=True
    close[spatula_22,pan_11]=True
    close[pan_11,spatula_22]=True
    on[knife_17,countertop_23]=True
    close[knife_17,countertop_23]=True
    close[countertop_23,knife_17]=True
    on[oil_9,countertop_23]=True
    close[oil_9,countertop_23]=True
    close[countertop_23,oil_9]=True
    on[sugar_10,countertop_23]=True
    close[sugar_10,countertop_23]=True
    close[countertop_23,sugar_10]=True
    on[salt_12,countertop_23]=True
    close[salt_12,countertop_23]=True
    close[countertop_23,salt_12]=True
    on[pepper_25,countertop_23]=True
    close[pepper_25,countertop_23]=True
    close[countertop_23,pepper_25]=True

    holds_lh[char,spatula_22]=True
    holds_rh[char,knife_17]=True


behavior prepare_tomato(tomato:item):
    body:
        achieve clean(tomato)        

behavior prepare_egg(egg:item, bowl:item):
    body:
        achieve inside(egg, bowl)
        achieve mixed(bowl)

behavior cook_scrambled_eggs_with_tomatoes(pan:item, stove:item, tomato:item, egg:item, sugar:item, salt:item, oil:item):
    body:
        achieve on(pan, stove)
        achieve is_on(stove)
        achieve inside(tomato, pan)
        achieve inside(egg, pan)
        achieve inside(sugar, pan)
        achieve inside(salt, pan)
        achieve inside(oil, pan)
        achieve mixed(pan)

behavior __goal__():
    body:
        bind pan: item where:
            is_pan(pan)
        bind stove: item where:
            is_stove(stove)
        bind tomato: item where:
            is_tomato(tomato)
        bind egg: item where:
            is_egg(egg)
        bind bowl: item where:
            is_bowl(bowl)
        bind sugar: item where:
            is_sugar(sugar)
        bind salt: item where:
            is_salt(salt)
        bind oil: item where:
            is_oil(oil)
        prepare_tomato(tomato)