Make spaghetti.
You can use a pot to process noodles. And process tomato, onion to make sause. Then mix them together to make spaghetti. However, I only have one pot and one pan.

behavior prepare_noodles(noodles:item, pot:item, stove:item):
    body:
        achieve boiled(noodles)

behavior prepare_sauce(tomato:item, onion:item, pan:item, stove:item):
    body:
        achieve sliced(tomato)
        achieve sliced(onion)
        achieve on(pan, stove)
        achieve is_on(stove)
        achieve inside(tomato, pan)
        achieve inside(onion, pan)
        achieve fried(tomato)
        achieve fried(onion)

behavior make_spaghetti(noodles:item, pot:item, stove:item, tomato:item, onion:item, pan:item):
    body:
        prepare_noodles(noodles, pot, stove)
        prepare_sauce(tomato, onion, pan, stove)
        bind countertop: item where:
            is_countertop(countertop)
        achieve on(pot, countertop)
        achieve on(pan, countertop)
        achieve inside(noodles, pan)
        achieve mixed(pan)
behavior __goal__():
    body:
        bind noodles: item where:
            is_noodles(noodles)
        bind pot: item where:
            is_pot(pot)
        bind tomato: item where:
            is_tomato(tomato)
        bind onion: item where:
            is_onion(onion)
        bind pan: item where:
            is_pan(pan)
        bind stove: item where:
            is_stove(stove)
        make_spaghetti(noodles, pot, stove, tomato, onion, pan)