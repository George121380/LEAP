problem "virtualhome-problem"
domain "virtualhome.cdl"

#!pragma planner_is_goal_serializable=False
#!pragma planner_is_goal_ordered=True
#!pragma planner_always_commit_skeleton=True

objects:
  basket:item
  char:character
  vegetables:item
  eggs:item
  cheese:item
  milk:item
  fridge:item

init:
  inside[vegetables,basket]=True
  inside[eggs,basket]=True
  inside[cheese,basket]=True
  inside[milk,basket]=True
  closed[fridge]=True
  closed[basket,fridge]=False

goal:
  is_off(light)


def all_foods_in_basket_in_fridge(basket: item):
  return inside[vegetables, fridge] and inside[eggs, fridge] and inside[cheese, fridge] and inside[milk, fridge] and closed[fridge]

behavior put_foods_in_fridge(basket: item):
  goal:
    all_foods_in_basket_in_fridge(basket)
  body:
    promotable:
      achieve inside(vegetables, basket)
      achieve inside(eggs, basket)
      achieve inside(cheese, basket)
      achieve inside(milk, basket)
      achieve closed(fridge)

goal:
  all_foods_in_basket_in_fridge(basket)

