problem "virtualhome-problem"
domain "virtualhome.cdl"

#!pragma planner_is_goal_serializable=False
#!pragma planner_is_goal_ordered=True
#!pragma planner_always_commit_skeleton=True

objects:
  bathroom_1:item
  floor_2:item
  floor_3:item
  floor_4:item
  floor_5:item
  floor_6:item
  floor_7:item
  floor_8:item
  wall_9:item
  wall_10:item
  wall_11:item
  wall_12:item
  wall_13:item
  wall_14:item
  ceiling_15:item
  ceiling_16:item
  ceiling_17:item
  ceiling_18:item
  ceiling_19:item
  ceiling_20:item
  mat_21:item
  curtain_22:item
  ceilinglamp_23:item
  walllamp_24:item
  walllamp_25:item
  walllamp_26:item
  bathroom_counter_27:item
  sink_28:item
  faucet_29:item
  bathtub_30:item
  towel_rack_31:item
  towel_rack_32:item
  towel_rack_33:item
  wallshelf_34:item
  shower_35:item
  bathroom_cabinet_36:item
  toilet_37:item
  shelf_38:item
  door_39:item
  doorjamb_40:item
  window_61:item
  light_62:item
  bedroom_64:item
  floor_65:item
  floor_66:item
  floor_67:item
  floor_68:item
  floor_69:item
  floor_70:item
  floor_71:item
  floor_72:item
  floor_73:item
  floor_74:item
  wall_75:item
  wall_76:item
  wall_77:item
  wall_78:item
  wall_79:item
  wall_80:item
  wall_81:item
  wall_82:item
  wall_83:item
  window_84:item
  ceiling_85:item
  ceiling_86:item
  ceiling_87:item
  ceiling_88:item
  ceiling_89:item
  ceiling_90:item
  ceiling_91:item
  ceiling_92:item
  ceiling_93:item
  ceilinglamp_94:item
  tablelamp_95:item
  chair_96:item
  bookshelf_97:item
  nightstand_98:item
  bed_99:item
  dresser_100:item
  chair_101:item
  hanger_102:item
  table_103:item
  doorjamb_104:item
  light_105:item
  mat_107:item
  drawing_108:item
  drawing_109:item
  drawing_110:item
  curtain_111:item
  curtain_112:item
  pillow_113:item
  pillow_114:item
  vase_115:item
  hanger_124:item
  hanger_125:item
  hanger_126:item
  hanger_127:item
  hanger_128:item
  hanger_129:item
  hanger_130:item
  hanger_131:item
  hanger_132:item
  hanger_133:item
  hanger_134:item
  closetdrawer_141:item
  closetdrawer_142:item
  closetdrawer_143:item
  closetdrawer_144:item
  closetdrawer_145:item
  closetdrawer_146:item
  dining_room_163:item
  floor_164:item
  floor_165:item
  floor_166:item
  floor_167:item
  floor_168:item
  floor_169:item
  floor_170:item
  wall_171:item
  wall_172:item
  wall_173:item
  wall_174:item
  wall_175:item
  wall_176:item
  ceiling_177:item
  ceiling_178:item
  ceiling_179:item
  ceiling_180:item
  ceiling_181:item
  ceiling_182:item
  door_183:item
  doorjamb_184:item
  maindoor_185:item
  ceilinglamp_186:item
  ceilinglamp_187:item
  tvstand_188:item
  table_189:item
  bench_190:item
  bench_191:item
  kitchen_counter_192:item
  sink_193:item
  faucet_194:item
  bookshelf_195:item
  mat_196:item
  drawing_197:item
  drawing_198:item
  orchid_199:item
  light_200:item
  powersocket_201:item
  television_202:item
  wall_clock_204:item
  phone_205:item
  photoframe_219:item
  cutting_board_223:item
  cutting_board_228:item
  oven_229:item
  tray_230:item
  toaster_231:item
  freezer_234:item
  stovefan_235:item
  coffe_maker_236:item
  microwave_238:item
  home_office_246:item
  floor_247:item
  floor_248:item
  floor_249:item
  floor_250:item
  floor_251:item
  floor_252:item
  floor_253:item
  floor_254:item
  floor_255:item
  wall_256:item
  wall_257:item
  wall_258:item
  wall_259:item
  wall_260:item
  wall_261:item
  wall_262:item
  wall_263:item
  ceiling_264:item
  ceiling_265:item
  ceiling_266:item
  ceiling_267:item
  ceiling_268:item
  ceiling_269:item
  ceiling_270:item
  ceiling_271:item
  ceiling_272:item
  doorjamb_273:item
  doorjamb_274:item
  window_275:item
  ceilinglamp_276:item
  walllamp_277:item
  walllamp_278:item
  couch_279:item
  bookshelf_280:item
  table_281:item
  desk_282:item
  chair_283:item
  dresser_284:item
  hanger_285:item
  hanger_287:item
  hanger_289:item
  hanger_291:item
  hanger_293:item
  hanger_295:item
  closetdrawer_296:item
  closetdrawer_299:item
  closetdrawer_301:item
  filing_cabinet_305:item
  standingmirror_306:item
  drawing_307:item
  mat_308:item
  drawing_309:item
  pillow_310:item
  curtain_311:item
  curtain_312:item
  curtain_313:item
  toy_314:item
  television_315:item
  light_316:item
  powersocket_317:item
  mouse_318:item
  mousepad_319:item
  cpuscreen_320:item
  computer_321:item
  keyboard_322:item
  cupboard_1000:item
  bowl_1001:item
  food_oatmeal_1002:item
  milk_1003:item
  ground_coffee_1004:item
  cup_1005:item
  juice_1006:item
  broom_2000:item
  knife_2001:item
  clothes_pants_2002:item
  blender_2003:item
  fork_2004:item
  piano_bench_2005:item
  pillow_2006:item
  shaving_cream_2007:item
  cup_2008:item
  food_food_2009:item
  clothes_skirt_2010:item
  towel_2011:item
  glue_2012:item
  food_jam_2013:item
  drawing_2014:item
  food_food_2015:item
  food_carrot_2016:item
  comb_2017:item
  stereo_2018:item
  food_food_2019:item
  band_aids_2020:item
  sheets_2021:item
  purse_2022:item
  laundry_detergent_2023:item
  food_food_2024:item
  clothes_shirt_2025:item
  check_2026:item
  mouthwash_2027:item
  video_game_controller_2028:item
  form_2029:item
  needle_2030:item
  button_2031:item
  wall_clock_2032:item
  rag_2033:item
  novel_2034:item
  fork_2035:item
  controller_2036:item
  centerpiece_2037:item
  food_rice_2038:item
  video_game_controller_2039:item
  clothes_pants_2040:item
  deck_of_cards_2041:item
  novel_2042:item
  juice_2043:item
  food_carrot_2044:item
  check_2045:item
  ground_coffee_2046:item
  piano_bench_2047:item
  blender_2048:item
  broom_2049:item
  pencil_2050:item
  check_2051:item
  food_food_2052:item
  oil_2053:item
  controller_2054:item
  food_food_2055:item
  stamp_2056:item
  food_salt_2057:item
  sheets_2058:item
  blow_dryer_2059:item
  check_2060:item
  bag_2061:item
  sheets_2062:item
  band_aids_2063:item
  char:character

init:
  clean[bathroom_1] = True
  is_room[bathroom_1]=True
  clean[floor_2] = True
  dirty[floor_3] = True
  dirty[floor_4] = True
  dirty[floor_5] = True
  dirty[floor_6] = True
  dirty[floor_7] = True
  clean[floor_8] = True
  dirty[wall_9] = True
  clean[wall_10] = True
  dirty[wall_11] = True
  dirty[wall_12] = True
  dirty[wall_13] = True
  dirty[wall_14] = True
  clean[ceiling_15] = True
  dirty[ceiling_16] = True
  dirty[ceiling_17] = True
  dirty[ceiling_18] = True
  clean[ceiling_19] = True
  clean[ceiling_20] = True
  dirty[mat_21] = True
  clean[curtain_22] = True
  closed[curtain_22] = True
  is_on[ceilinglamp_23] = True
  clean[ceilinglamp_23] = True
  is_on[walllamp_24] = True
  clean[walllamp_24] = True
  is_on[walllamp_25] = True
  clean[walllamp_25] = True
  is_on[walllamp_26] = True
  clean[walllamp_26] = True
  clean[bathroom_counter_27] = True
  closed[bathroom_counter_27] = True
  clean[sink_28] = True
  clean[faucet_29] = True
  is_off[faucet_29] = True
  clean[bathtub_30] = True
  clean[towel_rack_31] = True
  clean[towel_rack_32] = True
  clean[towel_rack_33] = True
  clean[wallshelf_34] = True
  clean[shower_35] = True
  clean[bathroom_cabinet_36] = True
  closed[bathroom_cabinet_36] = True
  closed[toilet_37] = True
  is_off[toilet_37] = True
  dirty[toilet_37] = True
  clean[shelf_38] = True
  clean[door_39] = True
  open[door_39] = True
  clean[doorjamb_40] = True
  open[doorjamb_40] = True
  clean[window_61] = True
  is_on[light_62] = True
  plugged[light_62] = True
  clean[light_62] = True
  clean[bedroom_64] = True
  is_room[bedroom_64]=True
  dirty[floor_65] = True
  clean[floor_66] = True
  clean[floor_67] = True
  clean[floor_68] = True
  clean[floor_69] = True
  dirty[floor_70] = True
  dirty[floor_71] = True
  dirty[floor_72] = True
  dirty[floor_73] = True
  dirty[floor_74] = True
  dirty[wall_75] = True
  clean[wall_76] = True
  clean[wall_77] = True
  clean[wall_78] = True
  clean[wall_79] = True
  dirty[wall_80] = True
  clean[wall_81] = True
  clean[wall_82] = True
  dirty[wall_83] = True
  clean[window_84] = True
  open[window_84] = True
  clean[ceiling_85] = True
  dirty[ceiling_86] = True
  clean[ceiling_87] = True
  clean[ceiling_88] = True
  clean[ceiling_89] = True
  dirty[ceiling_90] = True
  dirty[ceiling_91] = True
  clean[ceiling_92] = True
  dirty[ceiling_93] = True
  is_on[ceilinglamp_94] = True
  clean[ceilinglamp_94] = True
  is_on[tablelamp_95] = True
  clean[tablelamp_95] = True
  clean[chair_96] = True
  closed[bookshelf_97] = True
  dirty[bookshelf_97] = True
  clean[nightstand_98] = True
  open[nightstand_98] = True
  clean[bed_99] = True
  closed[dresser_100] = True
  dirty[dresser_100] = True
  clean[chair_101] = True
  clean[hanger_102] = True
  clean[table_103] = True
  clean[doorjamb_104] = True
  open[doorjamb_104] = True
  is_on[light_105] = True
  plugged[light_105] = True
  clean[light_105] = True
  dirty[mat_107] = True
  clean[drawing_108] = True
  clean[drawing_109] = True
  clean[drawing_110] = True
  clean[curtain_111] = True
  closed[curtain_111] = True
  clean[curtain_112] = True
  closed[curtain_112] = True
  clean[pillow_113] = True
  clean[pillow_114] = True
  clean[vase_115] = True
  clean[hanger_124] = True
  clean[hanger_125] = True
  clean[hanger_126] = True
  clean[hanger_127] = True
  clean[hanger_128] = True
  clean[hanger_129] = True
  clean[hanger_130] = True
  clean[hanger_131] = True
  clean[hanger_132] = True
  clean[hanger_133] = True
  clean[hanger_134] = True
  clean[closetdrawer_141] = True
  clean[closetdrawer_142] = True
  clean[closetdrawer_143] = True
  clean[closetdrawer_144] = True
  clean[closetdrawer_145] = True
  clean[closetdrawer_146] = True
  clean[dining_room_163] = True
  is_room[dining_room_163]=True
  clean[floor_164] = True
  dirty[floor_165] = True
  dirty[floor_166] = True
  dirty[floor_167] = True
  clean[floor_168] = True
  dirty[floor_169] = True
  clean[floor_170] = True
  dirty[wall_171] = True
  clean[wall_172] = True
  dirty[wall_173] = True
  clean[wall_174] = True
  clean[wall_175] = True
  dirty[wall_176] = True
  dirty[ceiling_177] = True
  dirty[ceiling_178] = True
  clean[ceiling_179] = True
  clean[ceiling_180] = True
  dirty[ceiling_181] = True
  dirty[ceiling_182] = True
  clean[door_183] = True
  open[door_183] = True
  clean[doorjamb_184] = True
  open[doorjamb_184] = True
  clean[maindoor_185] = True
  open[maindoor_185] = True
  is_on[ceilinglamp_186] = True
  clean[ceilinglamp_186] = True
  is_on[ceilinglamp_187] = True
  clean[ceilinglamp_187] = True
  clean[tvstand_188] = True
  clean[table_189] = True
  clean[bench_190] = True
  clean[bench_191] = True
  clean[kitchen_counter_192] = True
  closed[kitchen_counter_192] = True
  clean[sink_193] = True
  clean[faucet_194] = True
  is_off[faucet_194] = True
  clean[bookshelf_195] = True
  closed[bookshelf_195] = True
  clean[mat_196] = True
  clean[drawing_197] = True
  clean[drawing_198] = True
  clean[orchid_199] = True
  is_on[light_200] = True
  plugged[light_200] = True
  clean[light_200] = True
  clean[powersocket_201] = True
  is_on[television_202] = True
  plugged[television_202] = True
  clean[television_202] = True
  is_on[wall_clock_204] = True
  plugged[wall_clock_204] = True
  clean[wall_clock_204] = True
  clean[phone_205] = True
  is_off[phone_205] = True
  unplugged[phone_205] = True
  clean[photoframe_219] = True
  dirty[cutting_board_223] = True
  dirty[cutting_board_228] = True
  clean[oven_229] = True
  closed[oven_229] = True
  is_off[oven_229] = True
  plugged[oven_229] = True
  clean[tray_230] = True
  is_off[toaster_231] = True
  plugged[toaster_231] = True
  dirty[toaster_231] = True
  clean[freezer_234] = True
  closed[freezer_234] = True
  plugged[freezer_234] = True
  clean[stovefan_235] = True
  clean[coffe_maker_236] = True
  closed[coffe_maker_236] = True
  is_off[coffe_maker_236] = True
  plugged[coffe_maker_236] = True
  clean[microwave_238] = True
  closed[microwave_238] = True
  is_off[microwave_238] = True
  plugged[microwave_238] = True
  clean[home_office_246] = True
  is_room[home_office_246]=True
  dirty[floor_247] = True
  dirty[floor_248] = True
  dirty[floor_249] = True
  dirty[floor_250] = True
  clean[floor_251] = True
  dirty[floor_252] = True
  clean[floor_253] = True
  clean[floor_254] = True
  dirty[floor_255] = True
  dirty[wall_256] = True
  clean[wall_257] = True
  dirty[wall_258] = True
  dirty[wall_259] = True
  clean[wall_260] = True
  clean[wall_261] = True
  dirty[wall_262] = True
  dirty[wall_263] = True
  clean[ceiling_264] = True
  dirty[ceiling_265] = True
  clean[ceiling_266] = True
  clean[ceiling_267] = True
  clean[ceiling_268] = True
  clean[ceiling_269] = True
  dirty[ceiling_270] = True
  clean[ceiling_271] = True
  dirty[ceiling_272] = True
  clean[doorjamb_273] = True
  open[doorjamb_273] = True
  clean[doorjamb_274] = True
  open[doorjamb_274] = True
  clean[window_275] = True
  open[window_275] = True
  is_on[ceilinglamp_276] = True
  clean[ceilinglamp_276] = True
  is_on[walllamp_277] = True
  clean[walllamp_277] = True
  is_on[walllamp_278] = True
  clean[walllamp_278] = True
  dirty[couch_279] = True
  closed[bookshelf_280] = True
  dirty[bookshelf_280] = True
  clean[table_281] = True
  clean[desk_282] = True
  clean[chair_283] = True
  clean[dresser_284] = True
  closed[dresser_284] = True
  clean[hanger_285] = True
  clean[hanger_287] = True
  clean[hanger_289] = True
  clean[hanger_291] = True
  clean[hanger_293] = True
  clean[hanger_295] = True
  clean[closetdrawer_296] = True
  clean[closetdrawer_299] = True
  clean[closetdrawer_301] = True
  clean[filing_cabinet_305] = True
  closed[filing_cabinet_305] = True
  clean[standingmirror_306] = True
  clean[drawing_307] = True
  clean[mat_308] = True
  clean[drawing_309] = True
  clean[pillow_310] = True
  closed[curtain_311] = True
  dirty[curtain_311] = True
  clean[curtain_312] = True
  closed[curtain_312] = True
  closed[curtain_313] = True
  dirty[curtain_313] = True
  dirty[toy_314] = True
  clean[television_315] = True
  is_off[television_315] = True
  plugged[television_315] = True
  is_on[light_316] = True
  plugged[light_316] = True
  clean[light_316] = True
  clean[powersocket_317] = True
  clean[mouse_318] = True
  plugged[mouse_318] = True
  dirty[mousepad_319] = True
  clean[cpuscreen_320] = True
  is_on[computer_321] = True
  clean[computer_321] = True
  clean[keyboard_322] = True
  plugged[keyboard_322] = True
  clean[cupboard_1000] = True
  closed[cupboard_1000] = True
  clean[bowl_1001] = True
  clean[food_oatmeal_1002] = True
  clean[milk_1003] = True
  closed[milk_1003] = True
  clean[ground_coffee_1004] = True
  closed[ground_coffee_1004] = True
  clean[cup_1005] = True
  clean[juice_1006] = True
  clean[broom_2000] = True
  clean[knife_2001] = True
  clean[clothes_pants_2002] = True
  is_on[blender_2003] = True
  closed[blender_2003] = True
  plugged[blender_2003] = True
  clean[blender_2003] = True
  clean[fork_2004] = True
  clean[piano_bench_2005] = True
  clean[pillow_2006] = True
  clean[shaving_cream_2007] = True
  clean[cup_2008] = True
  dirty[food_food_2009] = True
  clean[clothes_skirt_2010] = True
  dirty[towel_2011] = True
  clean[glue_2012] = True
  clean[food_jam_2013] = True
  closed[food_jam_2013] = True
  clean[drawing_2014] = True
  clean[food_food_2015] = True
  dirty[food_carrot_2016] = True
  clean[comb_2017] = True
  clean[stereo_2018] = True
  closed[stereo_2018] = True
  unplugged[stereo_2018] = True
  clean[food_food_2019] = True
  clean[band_aids_2020] = True
  dirty[sheets_2021] = True
  clean[purse_2022] = True
  closed[purse_2022] = True
  clean[laundry_detergent_2023] = True
  dirty[food_food_2024] = True
  clean[clothes_shirt_2025] = True
  clean[check_2026] = True
  clean[mouthwash_2027] = True
  clean[video_game_controller_2028] = True
  is_off[video_game_controller_2028] = True
  plugged[video_game_controller_2028] = True
  clean[form_2029] = True
  clean[needle_2030] = True
  clean[button_2031] = True
  clean[wall_clock_2032] = True
  is_off[wall_clock_2032] = True
  plugged[wall_clock_2032] = True
  dirty[rag_2033] = True
  clean[novel_2034] = True
  closed[novel_2034] = True
  dirty[fork_2035] = True
  clean[controller_2036] = True
  plugged[controller_2036] = True
  clean[centerpiece_2037] = True
  clean[food_rice_2038] = True
  clean[video_game_controller_2039] = True
  unplugged[video_game_controller_2039] = True
  clean[clothes_pants_2040] = True
  clean[deck_of_cards_2041] = True
  clean[novel_2042] = True
  open[novel_2042] = True
  clean[juice_2043] = True
  dirty[food_carrot_2044] = True
  clean[check_2045] = True
  clean[ground_coffee_2046] = True
  closed[ground_coffee_2046] = True
  dirty[piano_bench_2047] = True
  clean[blender_2048] = True
  plugged[blender_2048] = True
  open[blender_2048] = True
  clean[broom_2049] = True
  clean[pencil_2050] = True
  clean[check_2051] = True
  dirty[food_food_2052] = True
  clean[oil_2053] = True
  clean[controller_2054] = True
  plugged[controller_2054] = True
  clean[food_food_2055] = True
  clean[stamp_2056] = True
  clean[food_salt_2057] = True
  clean[sheets_2058] = True
  clean[blow_dryer_2059] = True
  is_off[blow_dryer_2059] = True
  plugged[blow_dryer_2059] = True
  clean[check_2060] = True
  clean[bag_2061] = True
  open[bag_2061] = True
  clean[sheets_2062] = True
  clean[band_aids_2063] = True
  close[laundry_detergent_2023,filing_cabinet_305]=True
  close[food_rice_2038,kitchen_counter_192]=True
  facing[mat_107,drawing_109]=True
  facing[mat_107,drawing_110]=True
  close[video_game_controller_2028,table_103]=True
  close[juice_2043,freezer_234]=True
  inside[wall_80,bedroom_64]=True
  inside[deck_of_cards_2041,bedroom_64]=True
  inside[deck_of_cards_2041,dresser_100]=True
  on[cutting_board_228,microwave_238]=True
  close[doorjamb_273,hanger_128]=True
  close[doorjamb_273,hanger_129]=True
  close[doorjamb_273,wall_258]=True
  close[doorjamb_273,wall_257]=True
  close[doorjamb_273,wall_259]=True
  close[doorjamb_273,wall_11]=True
  close[doorjamb_273,ceiling_269]=True
  close[doorjamb_273,bookshelf_280]=True
  close[doorjamb_273,desk_282]=True
  close[doorjamb_273,shower_35]=True
  close[doorjamb_273,light_316]=True
  close[doorjamb_273,powersocket_317]=True
  close[doorjamb_273,mouse_318]=True
  close[doorjamb_273,mousepad_319]=True
  close[doorjamb_273,floor_72]=True
  close[doorjamb_273,wall_75]=True
  close[doorjamb_273,wall_82]=True
  close[doorjamb_273,wall_83]=True
  close[doorjamb_273,ceiling_91]=True
  close[doorjamb_273,chair_96]=True
  close[doorjamb_273,floor_252]=True
  close[doorjamb_273,hanger_125]=True
  on[table_103,floor_70]=True
  inside[piano_bench_2005,home_office_246]=True
  close[curtain_313,wall_256]=True
  close[curtain_313,wall_260]=True
  close[curtain_313,ceiling_266]=True
  close[curtain_313,ceiling_267]=True
  close[curtain_313,standingmirror_306]=True
  close[curtain_313,window_275]=True
  close[curtain_313,curtain_311]=True
  close[curtain_313,curtain_312]=True
  close[curtain_313,floor_250]=True
  close[curtain_313,couch_279]=True
  facing[ceilinglamp_186,drawing_197]=True
  facing[ceilinglamp_186,drawing_198]=True
  on[ceiling_180,wall_175]=True
  close[mousepad_319,hanger_128]=True
  close[mousepad_319,wall_257]=True
  close[mousepad_319,hanger_129]=True
  close[mousepad_319,hanger_130]=True
  close[mousepad_319,hanger_131]=True
  close[mousepad_319,wall_258]=True
  close[mousepad_319,closetdrawer_141]=True
  close[mousepad_319,closetdrawer_142]=True
  close[mousepad_319,closetdrawer_143]=True
  close[mousepad_319,closetdrawer_144]=True
  close[mousepad_319,doorjamb_273]=True
  close[mousepad_319,closetdrawer_146]=True
  close[mousepad_319,closetdrawer_145]=True
  close[mousepad_319,desk_282]=True
  close[mousepad_319,chair_283]=True
  close[mousepad_319,light_316]=True
  close[mousepad_319,powersocket_317]=True
  close[mousepad_319,mouse_318]=True
  close[mousepad_319,cpuscreen_320]=True
  close[mousepad_319,computer_321]=True
  close[mousepad_319,keyboard_322]=True
  close[mousepad_319,floor_71]=True
  close[mousepad_319,floor_72]=True
  close[mousepad_319,wall_75]=True
  close[mousepad_319,wall_83]=True
  close[mousepad_319,dresser_100]=True
  close[mousepad_319,floor_253]=True
  close[mousepad_319,floor_252]=True
  close[mousepad_319,hanger_125]=True
  close[mousepad_319,hanger_126]=True
  close[mousepad_319,hanger_127]=True
  on[food_food_2024,table_281]=True
  inside[food_food_2015,freezer_234]=True
  inside[food_food_2015,dining_room_163]=True
  close[curtain_22,towel_rack_32]=True
  close[curtain_22,wall_9]=True
  close[curtain_22,wall_10]=True
  close[curtain_22,wall_13]=True
  close[curtain_22,ceiling_18]=True
  close[curtain_22,ceiling_19]=True
  close[curtain_22,ceiling_20]=True
  close[curtain_22,window_61]=True
  close[curtain_22,bathtub_30]=True
  inside[sink_28,bathroom_1]=True
  inside[sink_28,bathroom_counter_27]=True
  facing[microwave_238,wall_clock_204]=True
  close[bathroom_counter_27,floor_2]=True
  close[bathroom_counter_27,floor_3]=True
  close[bathroom_counter_27,floor_4]=True
  close[bathroom_counter_27,wall_9]=True
  close[bathroom_counter_27,blow_dryer_2059]=True
  close[bathroom_counter_27,wall_12]=True
  close[bathroom_counter_27,mat_21]=True
  close[bathroom_counter_27,walllamp_24]=True
  close[bathroom_counter_27,walllamp_25]=True
  close[bathroom_counter_27,sink_28]=True
  close[bathroom_counter_27,faucet_29]=True
  close[bathroom_counter_27,towel_rack_33]=True
  close[bathroom_counter_27,wallshelf_34]=True
  close[bathroom_counter_27,bathroom_cabinet_36]=True
  close[bathroom_counter_27,floor_166]=True
  close[bathroom_counter_27,floor_167]=True
  close[bathroom_counter_27,wall_174]=True
  close[bathroom_counter_27,wall_176]=True
  close[bathroom_counter_27,wall_clock_204]=True
  close[bathroom_counter_27,phone_205]=True
  close[bathroom_counter_27,shaving_cream_2007]=True
  close[bathroom_counter_27,comb_2017]=True
  close[bathroom_counter_27,band_aids_2020]=True
  close[bathroom_counter_27,oven_229]=True
  close[bathroom_counter_27,tray_230]=True
  close[bathroom_counter_27,stovefan_235]=True
  close[bathroom_counter_27,mouthwash_2027]=True
  close[bathroom_counter_27,wall_clock_2032]=True
  inside[hanger_125,bedroom_64]=True
  inside[hanger_125,dresser_100]=True
  facing[ceiling_264,drawing_307]=True
  facing[ceiling_264,drawing_309]=True
  inside[doorjamb_273,home_office_246]=True
  close[floor_70,bed_99]=True
  close[floor_70,floor_67]=True
  close[floor_70,floor_69]=True
  close[floor_70,table_103]=True
  close[floor_70,floor_71]=True
  close[floor_70,floor_73]=True
  close[floor_70,mat_107]=True
  close[floor_70,vase_115]=True
  inside[drawing_309,home_office_246]=True
  close[wall_75,hanger_128]=True
  close[wall_75,hanger_129]=True
  close[wall_75,hanger_130]=True
  close[wall_75,hanger_131]=True
  close[wall_75,hanger_132]=True
  close[wall_75,hanger_133]=True
  close[wall_75,hanger_134]=True
  close[wall_75,wall_257]=True
  close[wall_75,wall_258]=True
  close[wall_75,closetdrawer_141]=True
  close[wall_75,closetdrawer_142]=True
  close[wall_75,closetdrawer_143]=True
  close[wall_75,closetdrawer_144]=True
  close[wall_75,closetdrawer_145]=True
  close[wall_75,closetdrawer_146]=True
  close[wall_75,ceiling_270]=True
  close[wall_75,doorjamb_273]=True
  close[wall_75,desk_282]=True
  close[wall_75,chair_283]=True
  close[wall_75,light_316]=True
  close[wall_75,powersocket_317]=True
  close[wall_75,mouse_318]=True
  close[wall_75,mousepad_319]=True
  close[wall_75,cpuscreen_320]=True
  close[wall_75,computer_321]=True
  close[wall_75,keyboard_322]=True
  close[wall_75,floor_71]=True
  close[wall_75,wall_78]=True
  close[wall_75,wall_83]=True
  close[wall_75,ceiling_90]=True
  close[wall_75,dresser_100]=True
  close[wall_75,floor_253]=True
  close[wall_75,hanger_124]=True
  close[wall_75,hanger_125]=True
  close[wall_75,hanger_126]=True
  close[wall_75,hanger_127]=True
  inside[floor_73,bedroom_64]=True
  close[tablelamp_95,nightstand_98]=True
  close[tablelamp_95,bed_99]=True
  close[tablelamp_95,floor_68]=True
  close[tablelamp_95,floor_67]=True
  close[tablelamp_95,mat_107]=True
  close[tablelamp_95,wall_77]=True
  close[tablelamp_95,wall_79]=True
  close[tablelamp_95,curtain_112]=True
  close[tablelamp_95,pillow_113]=True
  close[tablelamp_95,curtain_111]=True
  close[tablelamp_95,pillow_114]=True
  close[tablelamp_95,window_84]=True
  close[dresser_100,hanger_128]=True
  close[dresser_100,hanger_129]=True
  close[dresser_100,hanger_130]=True
  close[dresser_100,hanger_131]=True
  close[dresser_100,hanger_132]=True
  close[dresser_100,hanger_133]=True
  close[dresser_100,hanger_134]=True
  close[dresser_100,wall_257]=True
  close[dresser_100,wall_258]=True
  close[dresser_100,closetdrawer_141]=True
  close[dresser_100,closetdrawer_142]=True
  close[dresser_100,closetdrawer_143]=True
  close[dresser_100,closetdrawer_144]=True
  close[dresser_100,closetdrawer_145]=True
  close[dresser_100,closetdrawer_146]=True
  close[dresser_100,ceiling_270]=True
  close[dresser_100,bag_2061]=True
  close[dresser_100,band_aids_2063]=True
  close[dresser_100,desk_282]=True
  close[dresser_100,deck_of_cards_2041]=True
  close[dresser_100,light_316]=True
  close[dresser_100,powersocket_317]=True
  close[dresser_100,mouse_318]=True
  close[dresser_100,mousepad_319]=True
  close[dresser_100,cpuscreen_320]=True
  close[dresser_100,computer_321]=True
  close[dresser_100,keyboard_322]=True
  close[dresser_100,floor_71]=True
  close[dresser_100,wall_75]=True
  close[dresser_100,wall_78]=True
  close[dresser_100,broom_2000]=True
  close[dresser_100,wall_83]=True
  close[dresser_100,ceiling_90]=True
  close[dresser_100,clothes_shirt_2025]=True
  close[dresser_100,clothes_pants_2040]=True
  close[dresser_100,floor_253]=True
  close[dresser_100,hanger_124]=True
  close[dresser_100,hanger_125]=True
  close[dresser_100,hanger_126]=True
  close[dresser_100,hanger_127]=True
  inside[cup_2008,dining_room_163]=True
  inside[wall_257,home_office_246]=True
  inside[food_carrot_2044,dining_room_163]=True
  inside[toilet_37,bathroom_1]=True
  inside[toilet_37,shower_35]=True
  facing[ceiling_270,computer_321]=True
  close[ceilinglamp_23,wall_9]=True
  close[ceilinglamp_23,wall_10]=True
  close[ceilinglamp_23,wall_11]=True
  close[ceilinglamp_23,wall_12]=True
  close[ceilinglamp_23,ceiling_15]=True
  close[ceilinglamp_23,ceiling_16]=True
  close[ceilinglamp_23,ceiling_17]=True
  close[ceilinglamp_23,ceiling_18]=True
  close[ceilinglamp_23,ceiling_19]=True
  close[ceilinglamp_23,ceiling_20]=True
  inside[mat_21,bathroom_1]=True
  inside[mouse_318,home_office_246]=True
  facing[wall_172,television_202]=True
  facing[wall_172,drawing_197]=True
  facing[wall_172,drawing_198]=True
  close[floor_65,floor_66]=True
  close[floor_65,floor_67]=True
  close[floor_65,bed_99]=True
  close[floor_65,chair_101]=True
  close[floor_65,floor_71]=True
  close[floor_65,mat_107]=True
  close[floor_65,drawing_109]=True
  close[floor_65,wall_78]=True
  close[floor_65,closetdrawer_142]=True
  close[floor_65,closetdrawer_141]=True
  close[floor_65,closetdrawer_145]=True
  close[floor_65,pillow_114]=True
  inside[ceiling_266,home_office_246]=True
  inside[ceiling_92,bedroom_64]=True
  close[ceiling_90,hanger_128]=True
  close[ceiling_90,hanger_129]=True
  close[ceiling_90,hanger_130]=True
  close[ceiling_90,hanger_131]=True
  close[ceiling_90,hanger_132]=True
  close[ceiling_90,hanger_133]=True
  close[ceiling_90,hanger_134]=True
  close[ceiling_90,wall_257]=True
  close[ceiling_90,ceiling_270]=True
  close[ceiling_90,light_316]=True
  close[ceiling_90,cpuscreen_320]=True
  close[ceiling_90,wall_75]=True
  close[ceiling_90,wall_78]=True
  close[ceiling_90,ceiling_85]=True
  close[ceiling_90,ceiling_89]=True
  close[ceiling_90,ceiling_91]=True
  close[ceiling_90,ceilinglamp_94]=True
  close[ceiling_90,dresser_100]=True
  close[ceiling_90,hanger_124]=True
  close[ceiling_90,hanger_125]=True
  close[ceiling_90,hanger_126]=True
  close[ceiling_90,hanger_127]=True
  inside[mouthwash_2027,bathroom_1]=True
  close[hanger_285,hanger_289]=True
  close[hanger_285,hanger_291]=True
  close[hanger_285,wall_260]=True
  close[hanger_285,hanger_293]=True
  close[hanger_285,wall_262]=True
  close[hanger_285,hanger_295]=True
  close[hanger_285,closetdrawer_296]=True
  close[hanger_285,ceiling_265]=True
  close[hanger_285,ceiling_266]=True
  close[hanger_285,closetdrawer_299]=True
  close[hanger_285,closetdrawer_301]=True
  close[hanger_285,drawing_307]=True
  close[hanger_285,dresser_284]=True
  close[hanger_285,hanger_287]=True
  inside[doorjamb_40,bathroom_1]=True
  on[vase_115,table_103]=True
  close[pillow_113,nightstand_98]=True
  close[pillow_113,floor_67]=True
  close[pillow_113,bed_99]=True
  close[pillow_113,floor_68]=True
  close[pillow_113,mat_107]=True
  close[pillow_113,wall_77]=True
  close[pillow_113,curtain_111]=True
  close[pillow_113,curtain_112]=True
  close[pillow_113,wall_79]=True
  close[pillow_113,pillow_114]=True
  close[pillow_113,window_84]=True
  close[pillow_113,tablelamp_95]=True
  close[light_200,floor_164]=True
  close[light_200,floor_165]=True
  close[light_200,floor_168]=True
  close[light_200,powersocket_201]=True
  close[light_200,wall_171]=True
  close[light_200,wall_173]=True
  close[light_200,ceiling_177]=True
  close[light_200,ceiling_178]=True
  close[light_200,doorjamb_184]=True
  close[light_200,maindoor_185]=True
  inside[wall_76,bedroom_64]=True
  close[light_316,hanger_128]=True
  close[light_316,hanger_129]=True
  close[light_316,wall_258]=True
  close[light_316,wall_257]=True
  close[light_316,ceiling_269]=True
  close[light_316,ceiling_270]=True
  close[light_316,closetdrawer_143]=True
  close[light_316,closetdrawer_144]=True
  close[light_316,doorjamb_273]=True
  close[light_316,closetdrawer_146]=True
  close[light_316,bookshelf_280]=True
  close[light_316,desk_282]=True
  close[light_316,powersocket_317]=True
  close[light_316,mouse_318]=True
  close[light_316,mousepad_319]=True
  close[light_316,cpuscreen_320]=True
  close[light_316,computer_321]=True
  close[light_316,floor_71]=True
  close[light_316,floor_72]=True
  close[light_316,wall_75]=True
  close[light_316,wall_83]=True
  close[light_316,ceiling_90]=True
  close[light_316,ceiling_91]=True
  close[light_316,chair_96]=True
  close[light_316,dresser_100]=True
  close[light_316,floor_253]=True
  close[light_316,floor_252]=True
  close[light_316,hanger_125]=True
  close[light_316,hanger_127]=True
  inside[towel_2011,dining_room_163]=True
  inside[floor_4,bathroom_1]=True
  on[keyboard_322,desk_282]=True
  inside[food_food_2052,freezer_234]=True
  inside[food_food_2052,dining_room_163]=True
  inside[walllamp_24,bathroom_1]=True
  inside[computer_321,home_office_246]=True
  on[glue_2012,desk_282]=True
  on[maindoor_185,floor_168]=True
  close[window_61,towel_rack_32]=True
  close[window_61,floor_5]=True
  close[window_61,wall_9]=True
  close[window_61,wall_10]=True
  close[window_61,wall_13]=True
  close[window_61,ceiling_19]=True
  close[window_61,curtain_22]=True
  close[window_61,bathtub_30]=True
  inside[hanger_285,dresser_284]=True
  inside[hanger_285,home_office_246]=True
  close[floor_66,floor_65]=True
  close[floor_66,floor_67]=True
  close[floor_66,bed_99]=True
  close[floor_66,chair_101]=True
  close[floor_66,floor_71]=True
  close[floor_66,mat_107]=True
  close[floor_66,drawing_109]=True
  close[floor_66,wall_78]=True
  close[floor_66,closetdrawer_142]=True
  close[floor_66,closetdrawer_141]=True
  close[floor_66,closetdrawer_145]=True
  close[floor_66,pillow_114]=True
  facing[doorjamb_104,television_202]=True
  facing[doorjamb_104,drawing_108]=True
  facing[doorjamb_104,drawing_197]=True
  facing[doorjamb_104,drawing_198]=True
  close[floor_165,kitchen_counter_192]=True
  close[floor_165,sink_193]=True
  close[floor_165,faucet_194]=True
  close[floor_165,floor_164]=True
  close[floor_165,floor_166]=True
  close[floor_165,toaster_231]=True
  close[floor_165,floor_168]=True
  close[floor_165,powersocket_201]=True
  close[floor_165,light_200]=True
  close[floor_165,freezer_234]=True
  close[floor_165,coffe_maker_236]=True
  close[floor_165,wall_173]=True
  close[floor_165,microwave_238]=True
  close[floor_165,wall_174]=True
  close[floor_165,table_189]=True
  close[floor_165,bench_191]=True
  inside[ceiling_85,bedroom_64]=True
  inside[kitchen_counter_192,dining_room_163]=True
  inside[band_aids_2020,bathroom_1]=True
  inside[ceiling_269,home_office_246]=True
  inside[towel_rack_33,bathroom_1]=True
  facing[drawing_110,drawing_108]=True
  inside[floor_253,home_office_246]=True
  close[floor_3,floor_2]=True
  close[floor_3,floor_4]=True
  close[floor_3,floor_6]=True
  close[floor_3,wall_9]=True
  close[floor_3,wall_12]=True
  close[floor_3,mat_21]=True
  close[floor_3,walllamp_25]=True
  close[floor_3,bathroom_counter_27]=True
  close[floor_3,sink_28]=True
  close[floor_3,faucet_29]=True
  close[floor_3,towel_rack_31]=True
  close[floor_3,floor_167]=True
  close[floor_3,door_39]=True
  close[floor_3,wall_176]=True
  close[floor_3,door_183]=True
  close[floor_3,light_62]=True
  close[floor_3,floor_74]=True
  close[floor_3,phone_205]=True
  close[floor_3,wall_81]=True
  close[floor_3,oven_229]=True
  close[floor_3,tray_230]=True
  close[check_2051,filing_cabinet_305]=True
  close[floor_8,towel_rack_32]=True
  close[floor_8,floor_5]=True
  close[floor_8,shelf_38]=True
  close[floor_8,floor_7]=True
  close[floor_8,wall_10]=True
  close[floor_8,wall_11]=True
  close[floor_8,walllamp_26]=True
  close[floor_8,bathtub_30]=True
  close[stamp_2056,bookshelf_280]=True
  inside[floor_7,bathroom_1]=True
  on[bench_190,floor_168]=True
  inside[powersocket_201,dining_room_163]=True
  on[ceiling_20,wall_9]=True
  close[food_food_2015,freezer_234]=True
  close[needle_2030,filing_cabinet_305]=True
  close[band_aids_2020,bathroom_counter_27]=True
  inside[walllamp_278,home_office_246]=True
  close[fork_2035,cupboard_1000]=True
  inside[food_food_2055,dining_room_163]=True
  close[floor_167,floor_2]=True
  close[floor_167,floor_3]=True
  close[floor_167,wall_12]=True
  close[floor_167,mat_21]=True
  close[floor_167,walllamp_25]=True
  close[floor_167,bathroom_counter_27]=True
  close[floor_167,sink_28]=True
  close[floor_167,faucet_29]=True
  close[floor_167,floor_166]=True
  close[floor_167,floor_168]=True
  close[floor_167,floor_170]=True
  close[floor_167,wall_174]=True
  close[floor_167,wall_175]=True
  close[floor_167,wall_176]=True
  close[floor_167,door_183]=True
  close[floor_167,table_189]=True
  close[floor_167,bench_190]=True
  close[floor_167,bench_191]=True
  close[floor_167,mat_196]=True
  close[floor_167,orchid_199]=True
  close[floor_167,phone_205]=True
  close[floor_167,oven_229]=True
  close[floor_167,tray_230]=True
  close[wall_172,floor_168]=True
  close[wall_172,floor_169]=True
  close[wall_172,floor_170]=True
  close[wall_172,wall_171]=True
  close[wall_172,wall_175]=True
  close[wall_172,ceiling_178]=True
  close[wall_172,ceiling_179]=True
  close[wall_172,ceiling_180]=True
  close[wall_172,doorjamb_184]=True
  close[wall_172,maindoor_185]=True
  close[wall_172,ceilinglamp_186]=True
  close[wall_172,tvstand_188]=True
  close[wall_172,table_189]=True
  close[wall_172,bench_190]=True
  close[wall_172,bookshelf_195]=True
  close[wall_172,mat_196]=True
  close[wall_172,drawing_197]=True
  close[wall_172,orchid_199]=True
  close[wall_172,television_202]=True
  close[wall_172,photoframe_219]=True
  close[wall_172,cutting_board_223]=True
  close[ceilinglamp_187,wall_173]=True
  close[ceilinglamp_187,wall_174]=True
  close[ceilinglamp_187,ceiling_177]=True
  close[ceilinglamp_187,ceiling_178]=True
  close[ceilinglamp_187,ceiling_181]=True
  close[ceilinglamp_187,ceiling_182]=True
  on[closetdrawer_142,closetdrawer_145]=True
  inside[maindoor_185,dining_room_163]=True
  close[ceiling_265,hanger_289]=True
  close[ceiling_265,hanger_291]=True
  close[ceiling_265,wall_259]=True
  close[ceiling_265,hanger_293]=True
  close[ceiling_265,wall_262]=True
  close[ceiling_265,wall_260]=True
  close[ceiling_265,ceiling_264]=True
  close[ceiling_265,ceiling_266]=True
  close[ceiling_265,ceiling_268]=True
  close[ceiling_265,drawing_307]=True
  close[ceiling_265,ceilinglamp_276]=True
  close[ceiling_265,walllamp_277]=True
  close[ceiling_265,drawing_309]=True
  close[ceiling_265,toy_314]=True
  close[ceiling_265,hanger_285]=True
  close[ceiling_265,hanger_287]=True
  close[hanger_125,hanger_128]=True
  close[hanger_125,hanger_129]=True
  close[hanger_125,hanger_130]=True
  close[hanger_125,hanger_131]=True
  close[hanger_125,hanger_132]=True
  close[hanger_125,hanger_133]=True
  close[hanger_125,hanger_134]=True
  close[hanger_125,wall_257]=True
  close[hanger_125,wall_258]=True
  close[hanger_125,closetdrawer_141]=True
  close[hanger_125,ceiling_270]=True
  close[hanger_125,closetdrawer_143]=True
  close[hanger_125,closetdrawer_144]=True
  close[hanger_125,doorjamb_273]=True
  close[hanger_125,ceiling_269]=True
  close[hanger_125,desk_282]=True
  close[hanger_125,light_316]=True
  close[hanger_125,mouse_318]=True
  close[hanger_125,mousepad_319]=True
  close[hanger_125,cpuscreen_320]=True
  close[hanger_125,keyboard_322]=True
  close[hanger_125,wall_75]=True
  close[hanger_125,wall_83]=True
  close[hanger_125,ceiling_90]=True
  close[hanger_125,ceiling_91]=True
  close[hanger_125,dresser_100]=True
  close[hanger_125,hanger_124]=True
  close[hanger_125,hanger_126]=True
  close[hanger_125,hanger_127]=True
  facing[ceiling_265,drawing_307]=True
  facing[ceiling_265,drawing_309]=True
  on[broom_2049,floor_164]=True
  inside[blender_2048,cupboard_1000]=True
  inside[blender_2048,dining_room_163]=True
  on[controller_2036,table_281]=True
  close[wall_14,floor_6]=True
  close[wall_14,door_39]=True
  close[wall_14,doorjamb_40]=True
  close[wall_14,light_105]=True
  close[wall_14,floor_73]=True
  close[wall_14,wall_11]=True
  close[wall_14,drawing_108]=True
  close[wall_14,wall_12]=True
  close[wall_14,wall_80]=True
  close[wall_14,ceiling_16]=True
  close[wall_14,wall_82]=True
  close[wall_14,wall_81]=True
  close[wall_14,ceiling_92]=True
  close[wall_14,light_62]=True
  close[wall_14,towel_rack_31]=True
  close[sheets_2062,filing_cabinet_305]=True
  facing[door_183,television_202]=True
  facing[door_183,drawing_108]=True
  facing[door_183,drawing_197]=True
  facing[door_183,drawing_198]=True
  close[light_62,floor_2]=True
  close[light_62,floor_3]=True
  close[light_62,floor_6]=True
  close[light_62,door_39]=True
  close[light_62,doorjamb_40]=True
  close[light_62,light_105]=True
  close[light_62,floor_73]=True
  close[light_62,floor_74]=True
  close[light_62,drawing_108]=True
  close[light_62,wall_12]=True
  close[light_62,wall_14]=True
  close[light_62,ceiling_15]=True
  close[light_62,wall_80]=True
  close[light_62,ceiling_16]=True
  close[light_62,wall_81]=True
  close[light_62,ceiling_92]=True
  close[light_62,ceiling_93]=True
  close[light_62,towel_rack_31]=True
  facing[bookshelf_195,television_202]=True
  facing[bookshelf_195,drawing_108]=True
  close[floor_67,floor_65]=True
  close[floor_67,nightstand_98]=True
  close[floor_67,bed_99]=True
  close[floor_67,floor_68]=True
  close[floor_67,floor_66]=True
  close[floor_67,floor_70]=True
  close[floor_67,table_103]=True
  close[floor_67,chair_101]=True
  close[floor_67,mat_107]=True
  close[floor_67,wall_77]=True
  close[floor_67,wall_78]=True
  close[floor_67,curtain_111]=True
  close[floor_67,curtain_112]=True
  close[floor_67,pillow_113]=True
  close[floor_67,pillow_114]=True
  close[floor_67,vase_115]=True
  close[floor_67,window_84]=True
  close[floor_67,wall_79]=True
  close[floor_67,tablelamp_95]=True
  on[form_2029,bookshelf_97]=True
  inside[floor_168,dining_room_163]=True
  close[rag_2033,towel_rack_32]=True
  on[comb_2017,bathroom_counter_27]=True
  inside[wall_clock_204,dining_room_163]=True
  facing[photoframe_219,drawing_197]=True
  close[ceiling_272,wall_261]=True
  close[ceiling_272,ceiling_267]=True
  close[ceiling_272,ceiling_271]=True
  close[ceiling_272,pillow_310]=True
  close[ceiling_272,curtain_311]=True
  close[ceiling_272,curtain_312]=True
  facing[ceiling_86,drawing_109]=True
  on[ceiling_264,wall_259]=True
  facing[wall_173,wall_clock_204]=True
  on[controller_2054,table_281]=True
  close[toaster_231,kitchen_counter_192]=True
  close[toaster_231,sink_193]=True
  close[toaster_231,faucet_194]=True
  close[toaster_231,floor_164]=True
  close[toaster_231,floor_165]=True
  close[toaster_231,coffe_maker_236]=True
  close[toaster_231,wall_173]=True
  close[toaster_231,ceiling_177]=True
  inside[food_oatmeal_1002,cupboard_1000]=True
  inside[food_oatmeal_1002,dining_room_163]=True
  close[floor_250,wall_256]=True
  close[floor_250,wall_260]=True
  close[floor_250,floor_249]=True
  close[floor_250,table_281]=True
  close[floor_250,wall_261]=True
  close[floor_250,floor_251]=True
  close[floor_250,standingmirror_306]=True
  close[floor_250,window_275]=True
  close[floor_250,mat_308]=True
  close[floor_250,curtain_311]=True
  close[floor_250,curtain_312]=True
  close[floor_250,curtain_313]=True
  close[floor_250,television_315]=True
  close[floor_250,couch_279]=True
  close[floor_250,floor_255]=True
  inside[floor_249,home_office_246]=True
  close[ceiling_15,bathroom_cabinet_36]=True
  close[ceiling_15,wall_9]=True
  close[ceiling_15,stovefan_235]=True
  close[ceiling_15,drawing_108]=True
  close[ceiling_15,wall_clock_204]=True
  close[ceiling_15,wall_12]=True
  close[ceiling_15,phone_205]=True
  close[ceiling_15,wall_176]=True
  close[ceiling_15,ceiling_16]=True
  close[ceiling_15,wall_81]=True
  close[ceiling_15,ceiling_93]=True
  close[ceiling_15,ceiling_181]=True
  close[ceiling_15,ceiling_20]=True
  close[ceiling_15,ceilinglamp_23]=True
  close[ceiling_15,walllamp_25]=True
  close[ceiling_15,faucet_29]=True
  close[ceiling_15,light_62]=True
  close[ceiling_15,towel_rack_31]=True
  close[band_aids_2063,dresser_100]=True
  inside[cutting_board_223,dining_room_163]=True
  on[purse_2022,couch_279]=True
  close[novel_2034,table_189]=True
  facing[cutting_board_228,wall_clock_204]=True
  close[walllamp_277,wall_259]=True
  close[walllamp_277,wall_262]=True
  close[walllamp_277,ceiling_264]=True
  close[walllamp_277,ceiling_265]=True
  close[walllamp_277,filing_cabinet_305]=True
  close[walllamp_277,drawing_307]=True
  close[walllamp_277,drawing_309]=True
  close[walllamp_277,toy_314]=True
  close[chair_283,cpuscreen_320]=True
  close[chair_283,wall_257]=True
  close[chair_283,keyboard_322]=True
  close[chair_283,computer_321]=True
  close[chair_283,wall_263]=True
  close[chair_283,wall_75]=True
  close[chair_283,ceiling_270]=True
  close[chair_283,mat_308]=True
  close[chair_283,walllamp_278]=True
  close[chair_283,floor_254]=True
  close[chair_283,desk_282]=True
  close[chair_283,floor_253]=True
  close[chair_283,mouse_318]=True
  close[chair_283,mousepad_319]=True
  on[toilet_37,floor_7]=True
  close[light_105,floor_6]=True
  close[light_105,door_39]=True
  close[light_105,doorjamb_40]=True
  close[light_105,floor_73]=True
  close[light_105,floor_72]=True
  close[light_105,wall_11]=True
  close[light_105,floor_7]=True
  close[light_105,wall_14]=True
  close[light_105,wall_80]=True
  close[light_105,ceiling_16]=True
  close[light_105,wall_82]=True
  close[light_105,ceiling_17]=True
  close[light_105,ceiling_91]=True
  close[light_105,ceiling_92]=True
  close[light_105,light_62]=True
  inside[wall_171,dining_room_163]=True
  close[hanger_126,hanger_128]=True
  close[hanger_126,hanger_129]=True
  close[hanger_126,hanger_130]=True
  close[hanger_126,hanger_131]=True
  close[hanger_126,hanger_132]=True
  close[hanger_126,hanger_133]=True
  close[hanger_126,hanger_134]=True
  close[hanger_126,wall_257]=True
  close[hanger_126,wall_258]=True
  close[hanger_126,closetdrawer_141]=True
  close[hanger_126,closetdrawer_142]=True
  close[hanger_126,closetdrawer_143]=True
  close[hanger_126,closetdrawer_144]=True
  close[hanger_126,ceiling_270]=True
  close[hanger_126,ceiling_269]=True
  close[hanger_126,desk_282]=True
  close[hanger_126,mouse_318]=True
  close[hanger_126,mousepad_319]=True
  close[hanger_126,cpuscreen_320]=True
  close[hanger_126,keyboard_322]=True
  close[hanger_126,wall_75]=True
  close[hanger_126,wall_78]=True
  close[hanger_126,wall_83]=True
  close[hanger_126,ceiling_90]=True
  close[hanger_126,ceiling_91]=True
  close[hanger_126,dresser_100]=True
  close[hanger_126,hanger_124]=True
  close[hanger_126,hanger_125]=True
  close[hanger_126,hanger_127]=True
  facing[floor_252,drawing_307]=True
  facing[floor_252,drawing_309]=True
  close[mat_308,wall_256]=True
  close[mat_308,wall_261]=True
  close[mat_308,wall_263]=True
  close[mat_308,floor_251]=True
  close[mat_308,chair_283]=True
  close[mat_308,doorjamb_274]=True
  close[mat_308,window_275]=True
  close[mat_308,pillow_310]=True
  close[mat_308,couch_279]=True
  close[mat_308,curtain_312]=True
  close[mat_308,table_281]=True
  close[mat_308,floor_250]=True
  close[mat_308,television_315]=True
  close[mat_308,curtain_311]=True
  close[mat_308,floor_254]=True
  close[mat_308,floor_255]=True
  close[wall_13,towel_rack_32]=True
  close[wall_13,towel_rack_33]=True
  close[wall_13,wallshelf_34]=True
  close[wall_13,floor_5]=True
  close[wall_13,wall_9]=True
  close[wall_13,wall_10]=True
  close[wall_13,ceiling_19]=True
  close[wall_13,curtain_22]=True
  close[wall_13,window_61]=True
  close[wall_13,bathtub_30]=True
  close[bag_2061,dresser_100]=True
  close[ceiling_18,towel_rack_32]=True
  close[ceiling_18,shelf_38]=True
  close[ceiling_18,wall_10]=True
  close[ceiling_18,wall_11]=True
  close[ceiling_18,ceiling_17]=True
  close[ceiling_18,ceiling_19]=True
  close[ceiling_18,curtain_22]=True
  close[ceiling_18,ceilinglamp_23]=True
  close[ceiling_18,walllamp_26]=True
  close[towel_rack_33,wallshelf_34]=True
  close[towel_rack_33,floor_4]=True
  close[towel_rack_33,wall_9]=True
  close[towel_rack_33,wall_13]=True
  close[towel_rack_33,wall_174]=True
  close[towel_rack_33,ceiling_20]=True
  close[towel_rack_33,walllamp_24]=True
  close[towel_rack_33,bathroom_counter_27]=True
  facing[wall_260,television_315]=True
  facing[wall_260,drawing_307]=True
  inside[curtain_313,home_office_246]=True
  inside[ceiling_180,dining_room_163]=True
  close[check_2045,bookshelf_195]=True
  close[couch_279,wall_256]=True
  close[couch_279,clothes_skirt_2010]=True
  close[couch_279,wall_261]=True
  close[couch_279,sheets_2021]=True
  close[couch_279,curtain_313]=True
  close[couch_279,wall_263]=True
  close[couch_279,purse_2022]=True
  close[couch_279,floor_251]=True
  close[couch_279,doorjamb_274]=True
  close[couch_279,window_275]=True
  close[couch_279,mat_308]=True
  close[couch_279,clothes_pants_2002]=True
  close[couch_279,pillow_310]=True
  close[couch_279,curtain_311]=True
  close[couch_279,curtain_312]=True
  close[couch_279,table_281]=True
  close[couch_279,floor_250]=True
  close[couch_279,television_315]=True
  close[couch_279,floor_254]=True
  close[couch_279,floor_255]=True
  close[dresser_284,hanger_289]=True
  close[dresser_284,hanger_291]=True
  close[dresser_284,wall_260]=True
  close[dresser_284,hanger_293]=True
  close[dresser_284,wall_262]=True
  close[dresser_284,hanger_295]=True
  close[dresser_284,closetdrawer_296]=True
  close[dresser_284,ceiling_266]=True
  close[dresser_284,closetdrawer_299]=True
  close[dresser_284,closetdrawer_301]=True
  close[dresser_284,standingmirror_306]=True
  close[dresser_284,drawing_307]=True
  close[dresser_284,floor_249]=True
  close[dresser_284,hanger_285]=True
  close[dresser_284,hanger_287]=True
  inside[table_103,bedroom_64]=True
  inside[hanger_128,bedroom_64]=True
  inside[hanger_128,dresser_100]=True
  on[bathtub_30,floor_8]=True
  close[curtain_112,nightstand_98]=True
  close[curtain_112,bed_99]=True
  close[curtain_112,floor_67]=True
  close[curtain_112,mat_107]=True
  close[curtain_112,wall_77]=True
  close[curtain_112,curtain_111]=True
  close[curtain_112,wall_79]=True
  close[curtain_112,pillow_113]=True
  close[curtain_112,pillow_114]=True
  close[curtain_112,window_84]=True
  close[curtain_112,ceiling_86]=True
  close[curtain_112,ceiling_87]=True
  close[curtain_112,tablelamp_95]=True
  on[piano_bench_2005,floor_254]=True
  inside[floor_164,dining_room_163]=True
  inside[food_rice_2038,dining_room_163]=True
  on[freezer_234,floor_166]=True
  on[microwave_238,kitchen_counter_192]=True
  facing[floor_67,drawing_109]=True
  on[bookshelf_97,floor_69]=True
  close[hanger_134,hanger_128]=True
  close[hanger_134,hanger_129]=True
  close[hanger_134,hanger_130]=True
  close[hanger_134,hanger_131]=True
  close[hanger_134,hanger_132]=True
  close[hanger_134,hanger_133]=True
  close[hanger_134,wall_257]=True
  close[hanger_134,closetdrawer_141]=True
  close[hanger_134,closetdrawer_142]=True
  close[hanger_134,closetdrawer_143]=True
  close[hanger_134,closetdrawer_144]=True
  close[hanger_134,ceiling_270]=True
  close[hanger_134,desk_282]=True
  close[hanger_134,cpuscreen_320]=True
  close[hanger_134,keyboard_322]=True
  close[hanger_134,wall_75]=True
  close[hanger_134,wall_78]=True
  close[hanger_134,ceiling_85]=True
  close[hanger_134,ceiling_90]=True
  close[hanger_134,dresser_100]=True
  close[hanger_134,hanger_124]=True
  close[hanger_134,hanger_125]=True
  close[hanger_134,hanger_126]=True
  close[hanger_134,hanger_127]=True
  inside[orchid_199,dining_room_163]=True
  inside[chair_96,bedroom_64]=True
  close[wall_174,floor_4]=True
  close[wall_174,wall_9]=True
  close[wall_174,ceiling_20]=True
  close[wall_174,mat_21]=True
  close[wall_174,walllamp_24]=True
  close[wall_174,bathroom_counter_27]=True
  close[wall_174,sink_28]=True
  close[wall_174,faucet_29]=True
  close[wall_174,towel_rack_33]=True
  close[wall_174,wallshelf_34]=True
  close[wall_174,bathroom_cabinet_36]=True
  close[wall_174,floor_165]=True
  close[wall_174,floor_166]=True
  close[wall_174,floor_167]=True
  close[wall_174,floor_164]=True
  close[wall_174,wall_173]=True
  close[wall_174,wall_176]=True
  close[wall_174,ceiling_177]=True
  close[wall_174,ceiling_181]=True
  close[wall_174,ceiling_182]=True
  close[wall_174,ceilinglamp_187]=True
  close[wall_174,table_189]=True
  close[wall_174,bench_191]=True
  close[wall_174,kitchen_counter_192]=True
  close[wall_174,sink_193]=True
  close[wall_174,faucet_194]=True
  close[wall_174,mat_196]=True
  close[wall_174,orchid_199]=True
  close[wall_174,wall_clock_204]=True
  close[wall_174,cutting_board_228]=True
  close[wall_174,oven_229]=True
  close[wall_174,tray_230]=True
  close[wall_174,freezer_234]=True
  close[wall_174,stovefan_235]=True
  close[wall_174,coffe_maker_236]=True
  close[wall_174,microwave_238]=True
  close[wall_77,nightstand_98]=True
  close[wall_77,bed_99]=True
  close[wall_77,floor_67]=True
  close[wall_77,chair_101]=True
  close[wall_77,mat_107]=True
  close[wall_77,wall_78]=True
  close[wall_77,curtain_111]=True
  close[wall_77,curtain_112]=True
  close[wall_77,pillow_113]=True
  close[wall_77,pillow_114]=True
  close[wall_77,wall_79]=True
  close[wall_77,window_84]=True
  close[wall_77,ceiling_86]=True
  close[wall_77,tablelamp_95]=True
  close[floor_164,kitchen_counter_192]=True
  close[floor_164,sink_193]=True
  close[floor_164,faucet_194]=True
  close[floor_164,broom_2049]=True
  close[floor_164,floor_165]=True
  close[floor_164,floor_166]=True
  close[floor_164,toaster_231]=True
  close[floor_164,floor_168]=True
  close[floor_164,powersocket_201]=True
  close[floor_164,light_200]=True
  close[floor_164,freezer_234]=True
  close[floor_164,coffe_maker_236]=True
  close[floor_164,wall_173]=True
  close[floor_164,microwave_238]=True
  close[floor_164,wall_174]=True
  close[floor_164,table_189]=True
  close[floor_164,bench_191]=True
  close[ceiling_179,drawing_197]=True
  close[ceiling_179,wall_172]=True
  close[ceiling_179,wall_175]=True
  close[ceiling_179,ceiling_178]=True
  close[ceiling_179,ceiling_180]=True
  close[ceiling_179,ceilinglamp_186]=True
  inside[piano_bench_2047,home_office_246]=True
  inside[bookshelf_280,home_office_246]=True
  facing[floor_170,drawing_197]=True
  facing[floor_170,drawing_198]=True
  inside[floor_70,bedroom_64]=True
  close[keyboard_322,hanger_128]=True
  close[keyboard_322,wall_257]=True
  close[keyboard_322,hanger_130]=True
  close[keyboard_322,hanger_131]=True
  close[keyboard_322,hanger_132]=True
  close[keyboard_322,hanger_133]=True
  close[keyboard_322,hanger_129]=True
  close[keyboard_322,hanger_134]=True
  close[keyboard_322,wall_258]=True
  close[keyboard_322,closetdrawer_141]=True
  close[keyboard_322,closetdrawer_142]=True
  close[keyboard_322,closetdrawer_143]=True
  close[keyboard_322,closetdrawer_144]=True
  close[keyboard_322,closetdrawer_145]=True
  close[keyboard_322,closetdrawer_146]=True
  close[keyboard_322,desk_282]=True
  close[keyboard_322,chair_283]=True
  close[keyboard_322,mouse_318]=True
  close[keyboard_322,mousepad_319]=True
  close[keyboard_322,cpuscreen_320]=True
  close[keyboard_322,computer_321]=True
  close[keyboard_322,floor_71]=True
  close[keyboard_322,wall_75]=True
  close[keyboard_322,wall_83]=True
  close[keyboard_322,dresser_100]=True
  close[keyboard_322,hanger_125]=True
  close[keyboard_322,hanger_124]=True
  close[keyboard_322,floor_253]=True
  close[keyboard_322,hanger_126]=True
  close[keyboard_322,hanger_127]=True
  inside[button_2031,home_office_246]=True
  inside[hanger_131,bedroom_64]=True
  inside[hanger_131,dresser_100]=True
  on[hanger_102,floor_68]=True
  inside[hanger_289,dresser_284]=True
  inside[hanger_289,home_office_246]=True
  inside[vase_115,bedroom_64]=True
  facing[ceiling_272,television_315]=True
  close[clothes_shirt_2025,dresser_100]=True
  inside[closetdrawer_299,dresser_284]=True
  inside[closetdrawer_299,home_office_246]=True
  inside[wall_79,bedroom_64]=True
  close[ceiling_177,faucet_194]=True
  close[ceiling_177,cutting_board_228]=True
  close[ceiling_177,toaster_231]=True
  close[ceiling_177,light_200]=True
  close[ceiling_177,coffe_maker_236]=True
  close[ceiling_177,wall_173]=True
  close[ceiling_177,microwave_238]=True
  close[ceiling_177,wall_174]=True
  close[ceiling_177,ceiling_178]=True
  close[ceiling_177,ceiling_182]=True
  close[ceiling_177,ceilinglamp_187]=True
  close[ceiling_264,wall_259]=True
  close[ceiling_264,shower_35]=True
  close[ceiling_264,ceiling_265]=True
  close[ceiling_264,wall_11]=True
  close[ceiling_264,toy_314]=True
  close[ceiling_264,ceiling_269]=True
  close[ceiling_264,ceiling_17]=True
  close[ceiling_264,walllamp_277]=True
  close[ceiling_264,drawing_309]=True
  close[ceiling_264,bookshelf_280]=True
  close[ceiling_264,walllamp_26]=True
  inside[bed_99,bedroom_64]=True
  close[drawing_198,bookshelf_195]=True
  close[drawing_198,doorjamb_104]=True
  close[drawing_198,wall_76]=True
  close[drawing_198,drawing_110]=True
  close[drawing_198,wall_175]=True
  close[drawing_198,wall_81]=True
  close[drawing_198,ceiling_180]=True
  close[drawing_198,door_183]=True
  close[drawing_198,ceiling_88]=True
  close[drawing_198,ceiling_93]=True
  close[drawing_198,cutting_board_223]=True
  on[orchid_199,table_189]=True
  close[hanger_124,hanger_128]=True
  close[hanger_124,hanger_129]=True
  close[hanger_124,hanger_130]=True
  close[hanger_124,hanger_131]=True
  close[hanger_124,hanger_132]=True
  close[hanger_124,hanger_133]=True
  close[hanger_124,hanger_134]=True
  close[hanger_124,wall_257]=True
  close[hanger_124,wall_258]=True
  close[hanger_124,closetdrawer_141]=True
  close[hanger_124,closetdrawer_142]=True
  close[hanger_124,closetdrawer_143]=True
  close[hanger_124,closetdrawer_144]=True
  close[hanger_124,ceiling_270]=True
  close[hanger_124,ceiling_269]=True
  close[hanger_124,desk_282]=True
  close[hanger_124,cpuscreen_320]=True
  close[hanger_124,keyboard_322]=True
  close[hanger_124,wall_75]=True
  close[hanger_124,wall_78]=True
  close[hanger_124,wall_83]=True
  close[hanger_124,ceiling_85]=True
  close[hanger_124,ceiling_90]=True
  close[hanger_124,ceiling_91]=True
  close[hanger_124,dresser_100]=True
  close[hanger_124,hanger_125]=True
  close[hanger_124,hanger_126]=True
  close[hanger_124,hanger_127]=True
  inside[wall_263,home_office_246]=True
  close[television_202,drawing_197]=True
  close[television_202,floor_169]=True
  close[television_202,wall_171]=True
  close[television_202,wall_172]=True
  close[television_202,photoframe_219]=True
  close[television_202,tvstand_188]=True
  inside[drawing_2014,filing_cabinet_305]=True
  inside[drawing_2014,home_office_246]=True
  close[cutting_board_223,bookshelf_195]=True
  close[cutting_board_223,drawing_198]=True
  close[cutting_board_223,floor_169]=True
  close[cutting_board_223,floor_170]=True
  close[cutting_board_223,wall_172]=True
  close[cutting_board_223,wall_175]=True
  close[cutting_board_223,food_carrot_2044]=True
  close[microwave_238,kitchen_counter_192]=True
  close[microwave_238,sink_193]=True
  close[microwave_238,faucet_194]=True
  close[microwave_238,cutting_board_228]=True
  close[microwave_238,oven_229]=True
  close[microwave_238,floor_166]=True
  close[microwave_238,floor_165]=True
  close[microwave_238,floor_164]=True
  close[microwave_238,freezer_234]=True
  close[microwave_238,coffe_maker_236]=True
  close[microwave_238,wall_173]=True
  close[microwave_238,wall_174]=True
  close[microwave_238,ceiling_177]=True
  close[microwave_238,ceiling_182]=True
  inside[novel_2034,dining_room_163]=True
  facing[walllamp_278,computer_321]=True
  on[pencil_2050,table_103]=True
  on[filing_cabinet_305,floor_248]=True
  facing[oven_229,wall_clock_204]=True
  inside[wall_11,bathroom_1]=True
  inside[mat_308,home_office_246]=True
  inside[blow_dryer_2059,bathroom_1]=True
  facing[floor_253,computer_321]=True
  close[hanger_130,hanger_128]=True
  close[hanger_130,hanger_129]=True
  close[hanger_130,wall_257]=True
  close[hanger_130,hanger_131]=True
  close[hanger_130,hanger_132]=True
  close[hanger_130,hanger_133]=True
  close[hanger_130,hanger_134]=True
  close[hanger_130,wall_258]=True
  close[hanger_130,closetdrawer_141]=True
  close[hanger_130,closetdrawer_142]=True
  close[hanger_130,closetdrawer_143]=True
  close[hanger_130,closetdrawer_144]=True
  close[hanger_130,ceiling_270]=True
  close[hanger_130,ceiling_269]=True
  close[hanger_130,desk_282]=True
  close[hanger_130,mouse_318]=True
  close[hanger_130,mousepad_319]=True
  close[hanger_130,cpuscreen_320]=True
  close[hanger_130,keyboard_322]=True
  close[hanger_130,wall_75]=True
  close[hanger_130,wall_83]=True
  close[hanger_130,ceiling_90]=True
  close[hanger_130,ceiling_91]=True
  close[hanger_130,dresser_100]=True
  close[hanger_130,hanger_124]=True
  close[hanger_130,hanger_125]=True
  close[hanger_130,hanger_126]=True
  close[hanger_130,hanger_127]=True
  facing[ceiling_271,computer_321]=True
  facing[ceiling_271,television_315]=True
  close[knife_2001,table_281]=True
  close[sheets_2021,couch_279]=True
  close[milk_1003,freezer_234]=True
  on[ceiling_85,wall_78]=True
  inside[wall_256,home_office_246]=True
  close[check_2026,filing_cabinet_305]=True
  inside[wall_82,bedroom_64]=True
  close[wall_clock_2032,bathroom_counter_27]=True
  on[stereo_2018,table_103]=True
  inside[juice_2043,freezer_234]=True
  inside[juice_2043,dining_room_163]=True
  facing[wall_174,wall_clock_204]=True
  facing[wall_261,television_315]=True
  inside[shaving_cream_2007,bathroom_1]=True
  inside[floor_66,bedroom_64]=True
  inside[ceiling_20,bathroom_1]=True
  inside[knife_2001,home_office_246]=True
  close[floor_5,towel_rack_32]=True
  close[floor_5,floor_4]=True
  close[floor_5,floor_6]=True
  close[floor_5,floor_8]=True
  close[floor_5,wall_9]=True
  close[floor_5,wall_10]=True
  close[floor_5,wall_13]=True
  close[floor_5,mat_21]=True
  close[floor_5,window_61]=True
  close[floor_5,bathtub_30]=True
  close[oil_2053,table_189]=True
  inside[bathtub_30,bathroom_1]=True
  close[wall_10,towel_rack_32]=True
  close[wall_10,floor_5]=True
  close[wall_10,shelf_38]=True
  close[wall_10,floor_7]=True
  close[wall_10,floor_8]=True
  close[wall_10,wall_11]=True
  close[wall_10,wall_13]=True
  close[wall_10,ceiling_17]=True
  close[wall_10,ceiling_18]=True
  close[wall_10,ceiling_19]=True
  close[wall_10,curtain_22]=True
  close[wall_10,ceilinglamp_23]=True
  close[wall_10,walllamp_26]=True
  close[wall_10,window_61]=True
  close[wall_10,bathtub_30]=True
  close[walllamp_25,floor_2]=True
  close[walllamp_25,floor_3]=True
  close[walllamp_25,wall_12]=True
  close[walllamp_25,ceiling_15]=True
  close[walllamp_25,bathroom_counter_27]=True
  close[walllamp_25,towel_rack_31]=True
  close[walllamp_25,bathroom_cabinet_36]=True
  close[walllamp_25,floor_167]=True
  close[walllamp_25,floor_170]=True
  close[walllamp_25,wall_175]=True
  close[walllamp_25,wall_176]=True
  close[walllamp_25,ceiling_180]=True
  close[walllamp_25,ceiling_181]=True
  close[walllamp_25,door_183]=True
  close[walllamp_25,floor_74]=True
  close[walllamp_25,wall_clock_204]=True
  close[walllamp_25,phone_205]=True
  close[walllamp_25,wall_81]=True
  close[walllamp_25,ceiling_93]=True
  close[walllamp_25,doorjamb_104]=True
  close[walllamp_25,drawing_108]=True
  close[sheets_2058,bed_99]=True
  inside[hanger_127,bedroom_64]=True
  inside[hanger_127,dresser_100]=True
  facing[ceiling_88,drawing_108]=True
  facing[ceiling_88,drawing_110]=True
  inside[freezer_234,dining_room_163]=True
  close[centerpiece_2037,filing_cabinet_305]=True
  inside[curtain_311,curtain_312]=True
  inside[curtain_311,home_office_246]=True
  facing[curtain_112,drawing_109]=True
  close[ceiling_271,wall_257]=True
  close[ceiling_271,wall_261]=True
  close[ceiling_271,wall_263]=True
  close[ceiling_271,ceiling_268]=True
  close[ceiling_271,ceiling_270]=True
  close[ceiling_271,ceiling_272]=True
  close[ceiling_271,doorjamb_274]=True
  close[ceiling_271,ceilinglamp_276]=True
  close[ceiling_271,walllamp_278]=True
  inside[wall_75,bedroom_64]=True
  close[table_189,mat_196]=True
  close[table_189,floor_165]=True
  close[table_189,floor_166]=True
  close[table_189,floor_167]=True
  close[table_189,orchid_199]=True
  close[table_189,floor_168]=True
  close[table_189,floor_170]=True
  close[table_189,floor_169]=True
  close[table_189,floor_164]=True
  close[table_189,wall_172]=True
  close[table_189,wall_174]=True
  close[table_189,wall_173]=True
  close[table_189,wall_175]=True
  close[table_189,freezer_234]=True
  close[table_189,novel_2034]=True
  close[table_189,food_food_2055]=True
  close[table_189,video_game_controller_2039]=True
  close[table_189,oil_2053]=True
  close[table_189,bench_190]=True
  close[table_189,bench_191]=True
  close[ceilinglamp_276,ceiling_265]=True
  close[ceilinglamp_276,ceiling_267]=True
  close[ceilinglamp_276,ceiling_268]=True
  close[ceilinglamp_276,ceiling_269]=True
  close[ceilinglamp_276,ceiling_271]=True
  close[ceilinglamp_276,television_315]=True
  close[doorjamb_104,drawing_198]=True
  close[doorjamb_104,floor_74]=True
  close[doorjamb_104,floor_170]=True
  close[doorjamb_104,wall_76]=True
  close[doorjamb_104,phone_205]=True
  close[doorjamb_104,drawing_110]=True
  close[doorjamb_104,wall_175]=True
  close[doorjamb_104,wall_176]=True
  close[doorjamb_104,wall_81]=True
  close[doorjamb_104,wall_12]=True
  close[doorjamb_104,ceiling_180]=True
  close[doorjamb_104,door_183]=True
  close[doorjamb_104,walllamp_25]=True
  close[doorjamb_104,ceiling_93]=True
  facing[floor_66,drawing_109]=True
  inside[wall_259,home_office_246]=True
  inside[clothes_skirt_2010,home_office_246]=True
  facing[ceilinglamp_94,drawing_108]=True
  facing[ceilinglamp_94,drawing_109]=True
  facing[ceilinglamp_94,drawing_110]=True
  inside[door_39,bathroom_1]=True
  close[wall_12,floor_2]=True
  close[wall_12,floor_3]=True
  close[wall_12,floor_4]=True
  close[wall_12,floor_6]=True
  close[wall_12,wall_9]=True
  close[wall_12,wall_14]=True
  close[wall_12,ceiling_15]=True
  close[wall_12,ceiling_16]=True
  close[wall_12,ceiling_20]=True
  close[wall_12,mat_21]=True
  close[wall_12,ceilinglamp_23]=True
  close[wall_12,walllamp_25]=True
  close[wall_12,bathroom_counter_27]=True
  close[wall_12,sink_28]=True
  close[wall_12,faucet_29]=True
  close[wall_12,towel_rack_31]=True
  close[wall_12,bathroom_cabinet_36]=True
  close[wall_12,floor_167]=True
  close[wall_12,doorjamb_40]=True
  close[wall_12,door_39]=True
  close[wall_12,wall_176]=True
  close[wall_12,ceiling_181]=True
  close[wall_12,door_183]=True
  close[wall_12,light_62]=True
  close[wall_12,floor_74]=True
  close[wall_12,wall_clock_204]=True
  close[wall_12,phone_205]=True
  close[wall_12,wall_80]=True
  close[wall_12,wall_81]=True
  close[wall_12,ceiling_93]=True
  close[wall_12,oven_229]=True
  close[wall_12,tray_230]=True
  close[wall_12,doorjamb_104]=True
  close[wall_12,stovefan_235]=True
  close[wall_12,drawing_108]=True
  close[check_2060,filing_cabinet_305]=True
  inside[ceilinglamp_23,bathroom_1]=True
  close[towel_rack_32,floor_5]=True
  close[towel_rack_32,floor_8]=True
  close[towel_rack_32,wall_10]=True
  close[towel_rack_32,wall_13]=True
  close[towel_rack_32,rag_2033]=True
  close[towel_rack_32,ceiling_18]=True
  close[towel_rack_32,ceiling_19]=True
  close[towel_rack_32,curtain_22]=True
  close[towel_rack_32,window_61]=True
  close[towel_rack_32,bathtub_30]=True
  on[table_281,floor_251]=True
  close[hanger_131,hanger_128]=True
  close[hanger_131,hanger_129]=True
  close[hanger_131,hanger_130]=True
  close[hanger_131,wall_257]=True
  close[hanger_131,hanger_132]=True
  close[hanger_131,hanger_133]=True
  close[hanger_131,hanger_134]=True
  close[hanger_131,wall_258]=True
  close[hanger_131,closetdrawer_141]=True
  close[hanger_131,closetdrawer_142]=True
  close[hanger_131,closetdrawer_143]=True
  close[hanger_131,closetdrawer_144]=True
  close[hanger_131,ceiling_270]=True
  close[hanger_131,ceiling_269]=True
  close[hanger_131,desk_282]=True
  close[hanger_131,mouse_318]=True
  close[hanger_131,mousepad_319]=True
  close[hanger_131,cpuscreen_320]=True
  close[hanger_131,keyboard_322]=True
  close[hanger_131,wall_75]=True
  close[hanger_131,wall_83]=True
  close[hanger_131,ceiling_90]=True
  close[hanger_131,ceiling_91]=True
  close[hanger_131,dresser_100]=True
  close[hanger_131,hanger_124]=True
  close[hanger_131,hanger_125]=True
  close[hanger_131,hanger_126]=True
  close[hanger_131,hanger_127]=True
  facing[curtain_111,drawing_109]=True
  close[video_game_controller_2039,table_189]=True
  inside[ceiling_268,home_office_246]=True
  close[floor_69,bookshelf_97]=True
  close[floor_69,floor_68]=True
  close[floor_69,floor_70]=True
  close[floor_69,table_103]=True
  close[floor_69,floor_74]=True
  close[floor_69,mat_107]=True
  close[floor_69,wall_76]=True
  close[floor_69,drawing_110]=True
  close[floor_69,wall_79]=True
  close[floor_69,wall_81]=True
  close[floor_69,vase_115]=True
  close[floor_69,door_183]=True
  inside[ceilinglamp_94,bedroom_64]=True
  on[novel_2042,desk_282]=True
  close[food_carrot_2044,cutting_board_223]=True
  inside[form_2029,bedroom_64]=True
  close[vase_115,bed_99]=True
  close[vase_115,floor_67]=True
  close[vase_115,floor_69]=True
  close[vase_115,floor_70]=True
  close[vase_115,table_103]=True
  close[vase_115,mat_107]=True
  close[vase_115,wall_79]=True
  close[vase_115,ceiling_89]=True
  close[vase_115,ceilinglamp_94]=True
  inside[bench_191,dining_room_163]=True
  close[doorjamb_274,wall_257]=True
  close[doorjamb_274,wall_261]=True
  close[doorjamb_274,wall_263]=True
  close[doorjamb_274,ceiling_271]=True
  close[doorjamb_274,mat_308]=True
  close[doorjamb_274,walllamp_278]=True
  close[doorjamb_274,couch_279]=True
  close[doorjamb_274,floor_254]=True
  close[hanger_289,hanger_291]=True
  close[hanger_289,wall_260]=True
  close[hanger_289,hanger_293]=True
  close[hanger_289,wall_262]=True
  close[hanger_289,hanger_295]=True
  close[hanger_289,closetdrawer_296]=True
  close[hanger_289,ceiling_265]=True
  close[hanger_289,ceiling_266]=True
  close[hanger_289,closetdrawer_299]=True
  close[hanger_289,closetdrawer_301]=True
  close[hanger_289,drawing_307]=True
  close[hanger_289,dresser_284]=True
  close[hanger_289,hanger_285]=True
  close[hanger_289,hanger_287]=True
  close[hanger_295,hanger_289]=True
  close[hanger_295,hanger_291]=True
  close[hanger_295,wall_260]=True
  close[hanger_295,hanger_293]=True
  close[hanger_295,closetdrawer_296]=True
  close[hanger_295,ceiling_266]=True
  close[hanger_295,closetdrawer_299]=True
  close[hanger_295,closetdrawer_301]=True
  close[hanger_295,standingmirror_306]=True
  close[hanger_295,dresser_284]=True
  close[hanger_295,hanger_285]=True
  close[hanger_295,hanger_287]=True
  close[pillow_310,wall_261]=True
  close[pillow_310,ceiling_272]=True
  close[pillow_310,mat_308]=True
  close[pillow_310,couch_279]=True
  close[pillow_310,floor_255]=True
  inside[blender_2003,filing_cabinet_305]=True
  inside[blender_2003,home_office_246]=True
  facing[chair_101,drawing_109]=True
  close[toy_314,wall_259]=True
  close[toy_314,wall_262]=True
  close[toy_314,ceiling_264]=True
  close[toy_314,ceiling_265]=True
  close[toy_314,filing_cabinet_305]=True
  close[toy_314,drawing_307]=True
  close[toy_314,drawing_309]=True
  close[toy_314,walllamp_277]=True
  close[toy_314,floor_247]=True
  close[toy_314,floor_248]=True
  facing[doorjamb_273,drawing_309]=True
  inside[floor_6,bathroom_1]=True
  inside[controller_2054,home_office_246]=True
  inside[walllamp_26,bathroom_1]=True
  on[door_39,floor_73]=True
  on[door_39,floor_6]=True
  facing[floor_167,drawing_198]=True
  facing[floor_250,drawing_307]=True
  on[nightstand_98,mat_107]=True
  on[nightstand_98,floor_68]=True
  facing[ceiling_179,television_202]=True
  facing[ceiling_179,drawing_197]=True
  facing[ceiling_179,drawing_198]=True
  inside[hanger_287,dresser_284]=True
  inside[hanger_287,home_office_246]=True
  inside[doorjamb_184,dining_room_163]=True
  close[floor_71,wall_257]=True
  close[floor_71,closetdrawer_141]=True
  close[floor_71,closetdrawer_142]=True
  close[floor_71,closetdrawer_143]=True
  close[floor_71,closetdrawer_144]=True
  close[floor_71,closetdrawer_145]=True
  close[floor_71,closetdrawer_146]=True
  close[floor_71,desk_282]=True
  close[floor_71,light_316]=True
  close[floor_71,powersocket_317]=True
  close[floor_71,mouse_318]=True
  close[floor_71,mousepad_319]=True
  close[floor_71,cpuscreen_320]=True
  close[floor_71,computer_321]=True
  close[floor_71,keyboard_322]=True
  close[floor_71,floor_66]=True
  close[floor_71,floor_65]=True
  close[floor_71,floor_70]=True
  close[floor_71,floor_72]=True
  close[floor_71,wall_75]=True
  close[floor_71,wall_78]=True
  close[floor_71,dresser_100]=True
  close[floor_71,table_103]=True
  close[floor_71,mat_107]=True
  close[floor_71,floor_253]=True
  close[ceiling_86,wall_77]=True
  close[ceiling_86,wall_78]=True
  close[ceiling_86,curtain_111]=True
  close[ceiling_86,curtain_112]=True
  close[ceiling_86,wall_79]=True
  close[ceiling_86,window_84]=True
  close[ceiling_86,ceiling_85]=True
  close[ceiling_86,ceiling_87]=True
  close[ceiling_86,ceiling_89]=True
  close[ceiling_86,ceilinglamp_94]=True
  close[wall_76,bookshelf_97]=True
  close[wall_76,floor_69]=True
  close[wall_76,drawing_198]=True
  close[wall_76,doorjamb_104]=True
  close[wall_76,drawing_110]=True
  close[wall_76,wall_79]=True
  close[wall_76,wall_175]=True
  close[wall_76,wall_81]=True
  close[wall_76,door_183]=True
  close[wall_76,ceiling_88]=True
  close[ceiling_91,hanger_128]=True
  close[ceiling_91,hanger_129]=True
  close[ceiling_91,wall_258]=True
  close[ceiling_91,hanger_130]=True
  close[ceiling_91,hanger_131]=True
  close[ceiling_91,wall_11]=True
  close[ceiling_91,ceiling_269]=True
  close[ceiling_91,doorjamb_273]=True
  close[ceiling_91,ceiling_17]=True
  close[ceiling_91,shower_35]=True
  close[ceiling_91,light_316]=True
  close[ceiling_91,wall_82]=True
  close[ceiling_91,wall_83]=True
  close[ceiling_91,ceiling_90]=True
  close[ceiling_91,ceiling_92]=True
  close[ceiling_91,chair_96]=True
  close[ceiling_91,light_105]=True
  close[ceiling_91,hanger_124]=True
  close[ceiling_91,hanger_125]=True
  close[ceiling_91,hanger_126]=True
  close[ceiling_91,hanger_127]=True
  close[floor_169,bookshelf_195]=True
  close[floor_169,floor_168]=True
  close[floor_169,television_202]=True
  close[floor_169,floor_170]=True
  close[floor_169,wall_172]=True
  close[floor_169,wall_175]=True
  close[floor_169,photoframe_219]=True
  close[floor_169,tvstand_188]=True
  close[floor_169,table_189]=True
  close[floor_169,bench_190]=True
  close[floor_169,cutting_board_223]=True
  inside[faucet_194,dining_room_163]=True
  close[curtain_111,nightstand_98]=True
  close[curtain_111,bed_99]=True
  close[curtain_111,floor_67]=True
  close[curtain_111,mat_107]=True
  close[curtain_111,wall_77]=True
  close[curtain_111,wall_79]=True
  close[curtain_111,curtain_112]=True
  close[curtain_111,pillow_113]=True
  close[curtain_111,pillow_114]=True
  close[curtain_111,window_84]=True
  close[curtain_111,ceiling_86]=True
  close[curtain_111,ceiling_87]=True
  close[curtain_111,tablelamp_95]=True
  close[bench_190,mat_196]=True
  close[bench_190,floor_167]=True
  close[bench_190,floor_168]=True
  close[bench_190,orchid_199]=True
  close[bench_190,floor_170]=True
  close[bench_190,floor_169]=True
  close[bench_190,wall_172]=True
  close[bench_190,wall_175]=True
  close[bench_190,table_189]=True
  close[bench_190,bench_191]=True
  facing[floor_70,drawing_108]=True
  facing[floor_70,drawing_109]=True
  facing[floor_70,drawing_110]=True
  inside[shower_35,bathroom_1]=True
  inside[floor_255,home_office_246]=True
  facing[standingmirror_306,television_315]=True
  facing[standingmirror_306,drawing_307]=True
  on[shaving_cream_2007,bathroom_counter_27]=True
  close[hanger_128,hanger_129]=True
  close[hanger_128,hanger_130]=True
  close[hanger_128,hanger_131]=True
  close[hanger_128,hanger_132]=True
  close[hanger_128,hanger_133]=True
  close[hanger_128,hanger_134]=True
  close[hanger_128,wall_258]=True
  close[hanger_128,wall_257]=True
  close[hanger_128,closetdrawer_141]=True
  close[hanger_128,ceiling_270]=True
  close[hanger_128,closetdrawer_143]=True
  close[hanger_128,closetdrawer_144]=True
  close[hanger_128,doorjamb_273]=True
  close[hanger_128,ceiling_269]=True
  close[hanger_128,desk_282]=True
  close[hanger_128,light_316]=True
  close[hanger_128,mouse_318]=True
  close[hanger_128,mousepad_319]=True
  close[hanger_128,cpuscreen_320]=True
  close[hanger_128,keyboard_322]=True
  close[hanger_128,wall_75]=True
  close[hanger_128,wall_83]=True
  close[hanger_128,ceiling_90]=True
  close[hanger_128,ceiling_91]=True
  close[hanger_128,dresser_100]=True
  close[hanger_128,hanger_124]=True
  close[hanger_128,hanger_125]=True
  close[hanger_128,hanger_126]=True
  close[hanger_128,hanger_127]=True
  close[food_food_2024,table_281]=True
  on[coffe_maker_236,kitchen_counter_192]=True
  inside[floor_167,dining_room_163]=True
  close[wall_176,floor_2]=True
  close[wall_176,floor_3]=True
  close[wall_176,wall_9]=True
  close[wall_176,wall_12]=True
  close[wall_176,ceiling_15]=True
  close[wall_176,mat_21]=True
  close[wall_176,walllamp_25]=True
  close[wall_176,bathroom_counter_27]=True
  close[wall_176,sink_28]=True
  close[wall_176,faucet_29]=True
  close[wall_176,bathroom_cabinet_36]=True
  close[wall_176,floor_167]=True
  close[wall_176,wall_174]=True
  close[wall_176,wall_175]=True
  close[wall_176,ceiling_181]=True
  close[wall_176,door_183]=True
  close[wall_176,wall_clock_204]=True
  close[wall_176,phone_205]=True
  close[wall_176,wall_81]=True
  close[wall_176,oven_229]=True
  close[wall_176,tray_230]=True
  close[wall_176,doorjamb_104]=True
  close[wall_176,stovefan_235]=True
  inside[bowl_1001,cupboard_1000]=True
  inside[bowl_1001,dining_room_163]=True
  inside[ceilinglamp_187,dining_room_163]=True
  facing[coffe_maker_236,wall_clock_204]=True
  close[pillow_114,floor_65]=True
  close[pillow_114,nightstand_98]=True
  close[pillow_114,floor_67]=True
  close[pillow_114,bed_99]=True
  close[pillow_114,floor_66]=True
  close[pillow_114,mat_107]=True
  close[pillow_114,wall_77]=True
  close[pillow_114,wall_78]=True
  close[pillow_114,curtain_111]=True
  close[pillow_114,curtain_112]=True
  close[pillow_114,pillow_113]=True
  close[pillow_114,wall_79]=True
  close[pillow_114,window_84]=True
  close[pillow_114,tablelamp_95]=True
  facing[floor_248,drawing_307]=True
  facing[floor_248,drawing_309]=True
  on[bed_99,mat_107]=True
  on[bed_99,floor_67]=True
  on[tvstand_188,floor_169]=True
  facing[ceiling_89,drawing_108]=True
  facing[ceiling_89,drawing_109]=True
  facing[ceiling_89,drawing_110]=True
  on[wall_clock_2032,bathroom_counter_27]=True
  inside[floor_2,bathroom_1]=True
  facing[pillow_113,drawing_109]=True
  inside[pencil_2050,bedroom_64]=True
  facing[ceiling_268,computer_321]=True
  facing[ceiling_268,drawing_307]=True
  facing[ceiling_268,drawing_309]=True
  on[ceiling_15,wall_12]=True
  inside[floor_170,dining_room_163]=True
  close[ceiling_181,bathroom_cabinet_36]=True
  close[ceiling_181,stovefan_235]=True
  close[ceiling_181,wall_clock_204]=True
  close[ceiling_181,phone_205]=True
  close[ceiling_181,wall_12]=True
  close[ceiling_181,ceiling_15]=True
  close[ceiling_181,wall_176]=True
  close[ceiling_181,wall_175]=True
  close[ceiling_181,ceiling_178]=True
  close[ceiling_181,wall_174]=True
  close[ceiling_181,ceiling_180]=True
  close[ceiling_181,ceiling_182]=True
  close[ceiling_181,walllamp_25]=True
  close[ceiling_181,ceilinglamp_186]=True
  close[ceiling_181,ceilinglamp_187]=True
  close[ceiling_181,faucet_29]=True
  inside[hanger_134,bedroom_64]=True
  inside[hanger_134,dresser_100]=True
  close[oven_229,floor_2]=True
  close[oven_229,floor_3]=True
  close[oven_229,floor_4]=True
  close[oven_229,wall_9]=True
  close[oven_229,wall_12]=True
  close[oven_229,mat_21]=True
  close[oven_229,walllamp_24]=True
  close[oven_229,bathroom_counter_27]=True
  close[oven_229,sink_28]=True
  close[oven_229,faucet_29]=True
  close[oven_229,bathroom_cabinet_36]=True
  close[oven_229,floor_166]=True
  close[oven_229,floor_167]=True
  close[oven_229,wall_174]=True
  close[oven_229,wall_176]=True
  close[oven_229,kitchen_counter_192]=True
  close[oven_229,food_food_2019]=True
  close[oven_229,cutting_board_228]=True
  close[oven_229,tray_230]=True
  close[oven_229,freezer_234]=True
  close[oven_229,stovefan_235]=True
  close[oven_229,microwave_238]=True
  inside[ground_coffee_1004,dining_room_163]=True
  close[stovefan_235,bathroom_cabinet_36]=True
  close[stovefan_235,oven_229]=True
  close[stovefan_235,tray_230]=True
  close[stovefan_235,wall_9]=True
  close[stovefan_235,freezer_234]=True
  close[stovefan_235,wall_clock_204]=True
  close[stovefan_235,wall_12]=True
  close[stovefan_235,wall_174]=True
  close[stovefan_235,ceiling_15]=True
  close[stovefan_235,wall_176]=True
  close[stovefan_235,ceiling_20]=True
  close[stovefan_235,ceiling_181]=True
  close[stovefan_235,ceiling_182]=True
  close[stovefan_235,walllamp_24]=True
  close[stovefan_235,bathroom_counter_27]=True
  close[stovefan_235,sink_28]=True
  close[stovefan_235,faucet_29]=True
  facing[door_39,drawing_110]=True
  close[floor_4,towel_rack_33]=True
  close[floor_4,wallshelf_34]=True
  close[floor_4,floor_2]=True
  close[floor_4,floor_3]=True
  close[floor_4,oven_229]=True
  close[floor_4,tray_230]=True
  close[floor_4,floor_166]=True
  close[floor_4,floor_5]=True
  close[floor_4,wall_9]=True
  close[floor_4,wall_12]=True
  close[floor_4,wall_174]=True
  close[floor_4,mat_21]=True
  close[floor_4,walllamp_24]=True
  close[floor_4,bathroom_counter_27]=True
  close[floor_4,sink_28]=True
  close[floor_4,faucet_29]=True
  on[doorjamb_40,floor_73]=True
  on[doorjamb_40,floor_6]=True
  close[ceiling_19,towel_rack_32]=True
  close[ceiling_19,wall_9]=True
  close[ceiling_19,wall_10]=True
  close[ceiling_19,wall_13]=True
  close[ceiling_19,ceiling_16]=True
  close[ceiling_19,ceiling_18]=True
  close[ceiling_19,ceiling_20]=True
  close[ceiling_19,curtain_22]=True
  close[ceiling_19,ceilinglamp_23]=True
  close[ceiling_19,window_61]=True
  on[button_2031,table_281]=True
  close[walllamp_24,towel_rack_33]=True
  close[walllamp_24,wallshelf_34]=True
  close[walllamp_24,floor_4]=True
  close[walllamp_24,oven_229]=True
  close[walllamp_24,tray_230]=True
  close[walllamp_24,bathroom_cabinet_36]=True
  close[walllamp_24,floor_166]=True
  close[walllamp_24,wall_9]=True
  close[walllamp_24,freezer_234]=True
  close[walllamp_24,stovefan_235]=True
  close[walllamp_24,wall_174]=True
  close[walllamp_24,ceiling_20]=True
  close[walllamp_24,ceiling_182]=True
  close[walllamp_24,bathroom_counter_27]=True
  close[food_food_2052,freezer_234]=True
  close[pillow_2006,bench_191]=True
  close[towel_2011,kitchen_counter_192]=True
  inside[keyboard_322,home_office_246]=True
  close[button_2031,table_281]=True
  close[controller_2036,table_281]=True
  facing[light_200,drawing_197]=True
  close[door_183,floor_2]=True
  close[door_183,floor_3]=True
  close[door_183,floor_69]=True
  close[door_183,drawing_198]=True
  close[door_183,floor_167]=True
  close[door_183,doorjamb_104]=True
  close[door_183,floor_170]=True
  close[door_183,floor_74]=True
  close[door_183,wall_76]=True
  close[door_183,phone_205]=True
  close[door_183,drawing_110]=True
  close[door_183,wall_175]=True
  close[door_183,wall_176]=True
  close[door_183,wall_81]=True
  close[door_183,wall_12]=True
  close[door_183,walllamp_25]=True
  close[wall_262,hanger_289]=True
  close[wall_262,hanger_291]=True
  close[wall_262,wall_259]=True
  close[wall_262,hanger_293]=True
  close[wall_262,wall_260]=True
  close[wall_262,closetdrawer_296]=True
  close[wall_262,ceiling_265]=True
  close[wall_262,closetdrawer_301]=True
  close[wall_262,filing_cabinet_305]=True
  close[wall_262,drawing_307]=True
  close[wall_262,walllamp_277]=True
  close[wall_262,drawing_309]=True
  close[wall_262,floor_248]=True
  close[wall_262,toy_314]=True
  close[wall_262,dresser_284]=True
  close[wall_262,hanger_285]=True
  close[wall_262,hanger_287]=True
  close[tvstand_188,drawing_197]=True
  close[tvstand_188,floor_168]=True
  close[tvstand_188,floor_169]=True
  close[tvstand_188,television_202]=True
  close[tvstand_188,wall_171]=True
  close[tvstand_188,wall_172]=True
  close[tvstand_188,photoframe_219]=True
  close[ceiling_266,hanger_289]=True
  close[ceiling_266,hanger_291]=True
  close[ceiling_266,wall_260]=True
  close[ceiling_266,hanger_293]=True
  close[ceiling_266,hanger_295]=True
  close[ceiling_266,ceiling_265]=True
  close[ceiling_266,ceiling_267]=True
  close[ceiling_266,standingmirror_306]=True
  close[ceiling_266,drawing_307]=True
  close[ceiling_266,curtain_313]=True
  close[ceiling_266,dresser_284]=True
  close[ceiling_266,hanger_285]=True
  close[ceiling_266,hanger_287]=True
  close[table_281,wall_261]=True
  close[table_281,controller_2054]=True
  close[table_281,food_food_2024]=True
  close[table_281,floor_251]=True
  close[table_281,button_2031]=True
  close[table_281,knife_2001]=True
  close[table_281,mat_308]=True
  close[table_281,controller_2036]=True
  close[table_281,couch_279]=True
  close[table_281,floor_248]=True
  close[table_281,floor_250]=True
  close[table_281,television_315]=True
  close[table_281,floor_254]=True
  close[table_281,floor_255]=True
  close[hanger_287,hanger_289]=True
  close[hanger_287,hanger_291]=True
  close[hanger_287,wall_260]=True
  close[hanger_287,hanger_293]=True
  close[hanger_287,wall_262]=True
  close[hanger_287,hanger_295]=True
  close[hanger_287,closetdrawer_296]=True
  close[hanger_287,ceiling_265]=True
  close[hanger_287,ceiling_266]=True
  close[hanger_287,closetdrawer_299]=True
  close[hanger_287,closetdrawer_301]=True
  close[hanger_287,standingmirror_306]=True
  close[hanger_287,dresser_284]=True
  close[hanger_287,hanger_285]=True
  inside[wall_173,dining_room_163]=True
  inside[ceiling_86,bedroom_64]=True
  facing[ceiling_178,television_202]=True
  facing[ceiling_178,drawing_197]=True
  facing[ceiling_178,drawing_198]=True
  on[ceiling_87,wall_79]=True
  inside[sheets_2021,home_office_246]=True
  on[band_aids_2020,bathroom_counter_27]=True
  on[cup_2008,kitchen_counter_192]=True
  close[shelf_38,floor_8]=True
  close[shelf_38,wall_10]=True
  close[shelf_38,ceiling_18]=True
  close[shelf_38,bathtub_30]=True
  on[desk_282,floor_253]=True
  facing[window_84,drawing_109]=True
  facing[wall_256,television_315]=True
  inside[light_105,bedroom_64]=True
  inside[television_315,home_office_246]=True
  close[wall_78,hanger_132]=True
  close[wall_78,hanger_133]=True
  close[wall_78,hanger_134]=True
  close[wall_78,closetdrawer_141]=True
  close[wall_78,closetdrawer_142]=True
  close[wall_78,closetdrawer_145]=True
  close[wall_78,floor_65]=True
  close[wall_78,floor_66]=True
  close[wall_78,floor_67]=True
  close[wall_78,floor_71]=True
  close[wall_78,wall_75]=True
  close[wall_78,wall_77]=True
  close[wall_78,window_84]=True
  close[wall_78,ceiling_85]=True
  close[wall_78,ceiling_86]=True
  close[wall_78,ceiling_90]=True
  close[wall_78,bed_99]=True
  close[wall_78,dresser_100]=True
  close[wall_78,chair_101]=True
  close[wall_78,mat_107]=True
  close[wall_78,drawing_109]=True
  close[wall_78,pillow_114]=True
  close[wall_78,hanger_124]=True
  close[wall_78,hanger_126]=True
  close[floor_68,bookshelf_97]=True
  close[floor_68,nightstand_98]=True
  close[floor_68,floor_67]=True
  close[floor_68,bed_99]=True
  close[floor_68,floor_69]=True
  close[floor_68,hanger_102]=True
  close[floor_68,mat_107]=True
  close[floor_68,wall_79]=True
  close[floor_68,pillow_113]=True
  close[floor_68,tablelamp_95]=True
  inside[ceiling_182,dining_room_163]=True
  close[wall_83,hanger_128]=True
  close[wall_83,hanger_129]=True
  close[wall_83,wall_258]=True
  close[wall_83,hanger_130]=True
  close[wall_83,hanger_131]=True
  close[wall_83,wall_259]=True
  close[wall_83,wall_257]=True
  close[wall_83,wall_11]=True
  close[wall_83,ceiling_269]=True
  close[wall_83,closetdrawer_143]=True
  close[wall_83,closetdrawer_144]=True
  close[wall_83,doorjamb_273]=True
  close[wall_83,closetdrawer_146]=True
  close[wall_83,bookshelf_280]=True
  close[wall_83,desk_282]=True
  close[wall_83,shower_35]=True
  close[wall_83,toilet_37]=True
  close[wall_83,light_316]=True
  close[wall_83,powersocket_317]=True
  close[wall_83,mouse_318]=True
  close[wall_83,mousepad_319]=True
  close[wall_83,cpuscreen_320]=True
  close[wall_83,computer_321]=True
  close[wall_83,keyboard_322]=True
  close[wall_83,floor_72]=True
  close[wall_83,wall_75]=True
  close[wall_83,wall_82]=True
  close[wall_83,ceiling_91]=True
  close[wall_83,chair_96]=True
  close[wall_83,dresser_100]=True
  close[wall_83,hanger_124]=True
  close[wall_83,floor_252]=True
  close[wall_83,hanger_125]=True
  close[wall_83,hanger_126]=True
  close[wall_83,hanger_127]=True
  facing[drawing_108,drawing_198]=True
  facing[drawing_108,drawing_110]=True
  close[cup_1005,freezer_234]=True
  on[knife_2001,table_281]=True
  inside[needle_2030,filing_cabinet_305]=True
  inside[needle_2030,home_office_246]=True
  inside[couch_279,home_office_246]=True
  inside[ceiling_89,bedroom_64]=True
  inside[hanger_130,bedroom_64]=True
  inside[hanger_130,dresser_100]=True
  inside[food_food_2024,home_office_246]=True
  close[floor_247,floor_248]=True
  close[floor_247,chair_96]=True
  close[floor_247,wall_259]=True
  close[floor_247,shower_35]=True
  close[floor_247,toilet_37]=True
  close[floor_247,floor_7]=True
  close[floor_247,wall_11]=True
  close[floor_247,toy_314]=True
  close[floor_247,filing_cabinet_305]=True
  close[floor_247,bookshelf_280]=True
  close[floor_247,walllamp_26]=True
  close[floor_247,floor_252]=True
  facing[floor_249,drawing_307]=True
  facing[couch_279,television_315]=True
  inside[nightstand_98,bedroom_64]=True
  close[wall_81,floor_2]=True
  close[wall_81,floor_3]=True
  close[wall_81,wall_12]=True
  close[wall_81,wall_14]=True
  close[wall_81,ceiling_15]=True
  close[wall_81,walllamp_25]=True
  close[wall_81,towel_rack_31]=True
  close[wall_81,door_39]=True
  close[wall_81,doorjamb_40]=True
  close[wall_81,floor_170]=True
  close[wall_81,wall_175]=True
  close[wall_81,wall_176]=True
  close[wall_81,ceiling_180]=True
  close[wall_81,door_183]=True
  close[wall_81,light_62]=True
  close[wall_81,floor_69]=True
  close[wall_81,drawing_198]=True
  close[wall_81,floor_73]=True
  close[wall_81,floor_74]=True
  close[wall_81,wall_76]=True
  close[wall_81,phone_205]=True
  close[wall_81,wall_80]=True
  close[wall_81,ceiling_88]=True
  close[wall_81,ceiling_92]=True
  close[wall_81,ceiling_93]=True
  close[wall_81,doorjamb_104]=True
  close[wall_81,drawing_108]=True
  close[wall_81,drawing_110]=True
  close[floor_168,mat_196]=True
  close[floor_168,floor_164]=True
  close[floor_168,floor_165]=True
  close[floor_168,orchid_199]=True
  close[floor_168,light_200]=True
  close[floor_168,powersocket_201]=True
  close[floor_168,floor_169]=True
  close[floor_168,wall_171]=True
  close[floor_168,floor_167]=True
  close[floor_168,wall_172]=True
  close[floor_168,wall_173]=True
  close[floor_168,doorjamb_184]=True
  close[floor_168,maindoor_185]=True
  close[floor_168,tvstand_188]=True
  close[floor_168,table_189]=True
  close[floor_168,bench_190]=True
  close[floor_168,bench_191]=True
  inside[desk_282,home_office_246]=True
  close[hanger_102,bookshelf_97]=True
  close[hanger_102,floor_68]=True
  close[hanger_102,ceiling_87]=True
  close[hanger_102,wall_79]=True
  inside[drawing_108,bedroom_64]=True
  facing[television_315,computer_321]=True
  facing[television_315,drawing_307]=True
  facing[television_315,drawing_309]=True
  inside[light_62,bathroom_1]=True
  inside[rag_2033,bathroom_1]=True
  close[hanger_127,hanger_128]=True
  close[hanger_127,hanger_129]=True
  close[hanger_127,hanger_130]=True
  close[hanger_127,hanger_131]=True
  close[hanger_127,hanger_132]=True
  close[hanger_127,hanger_133]=True
  close[hanger_127,hanger_134]=True
  close[hanger_127,wall_257]=True
  close[hanger_127,wall_258]=True
  close[hanger_127,closetdrawer_141]=True
  close[hanger_127,closetdrawer_142]=True
  close[hanger_127,closetdrawer_143]=True
  close[hanger_127,closetdrawer_144]=True
  close[hanger_127,ceiling_270]=True
  close[hanger_127,ceiling_269]=True
  close[hanger_127,desk_282]=True
  close[hanger_127,light_316]=True
  close[hanger_127,mouse_318]=True
  close[hanger_127,mousepad_319]=True
  close[hanger_127,cpuscreen_320]=True
  close[hanger_127,keyboard_322]=True
  close[hanger_127,wall_75]=True
  close[hanger_127,wall_83]=True
  close[hanger_127,ceiling_90]=True
  close[hanger_127,ceiling_91]=True
  close[hanger_127,dresser_100]=True
  close[hanger_127,hanger_124]=True
  close[hanger_127,hanger_125]=True
  close[hanger_127,hanger_126]=True
  close[closetdrawer_301,hanger_289]=True
  close[closetdrawer_301,hanger_291]=True
  close[closetdrawer_301,wall_260]=True
  close[closetdrawer_301,hanger_293]=True
  close[closetdrawer_301,wall_262]=True
  close[closetdrawer_301,hanger_295]=True
  close[closetdrawer_301,closetdrawer_296]=True
  close[closetdrawer_301,closetdrawer_299]=True
  close[closetdrawer_301,drawing_307]=True
  close[closetdrawer_301,floor_248]=True
  close[closetdrawer_301,floor_249]=True
  close[closetdrawer_301,dresser_284]=True
  close[closetdrawer_301,hanger_285]=True
  close[closetdrawer_301,hanger_287]=True
  facing[ceiling_269,drawing_307]=True
  facing[ceiling_269,drawing_309]=True
  inside[comb_2017,bathroom_1]=True
  on[food_carrot_2044,cutting_board_223]=True
  close[faucet_29,floor_2]=True
  close[faucet_29,floor_3]=True
  close[faucet_29,floor_4]=True
  close[faucet_29,wall_9]=True
  close[faucet_29,wall_12]=True
  close[faucet_29,ceiling_15]=True
  close[faucet_29,ceiling_20]=True
  close[faucet_29,mat_21]=True
  close[faucet_29,bathroom_counter_27]=True
  close[faucet_29,sink_28]=True
  close[faucet_29,bathroom_cabinet_36]=True
  close[faucet_29,floor_166]=True
  close[faucet_29,floor_167]=True
  close[faucet_29,wall_174]=True
  close[faucet_29,wall_176]=True
  close[faucet_29,ceiling_181]=True
  close[faucet_29,ceiling_182]=True
  close[faucet_29,wall_clock_204]=True
  close[faucet_29,oven_229]=True
  close[faucet_29,tray_230]=True
  close[faucet_29,stovefan_235]=True
  close[wallshelf_34,towel_rack_33]=True
  close[wallshelf_34,floor_4]=True
  close[wallshelf_34,wall_9]=True
  close[wallshelf_34,wall_13]=True
  close[wallshelf_34,wall_174]=True
  close[wallshelf_34,ceiling_20]=True
  close[wallshelf_34,walllamp_24]=True
  close[wallshelf_34,bathroom_counter_27]=True
  inside[floor_250,home_office_246]=True
  inside[hanger_291,dresser_284]=True
  inside[hanger_291,home_office_246]=True
  facing[orchid_199,drawing_197]=True
  facing[orchid_199,drawing_198]=True
  inside[closetdrawer_301,dresser_284]=True
  inside[closetdrawer_301,home_office_246]=True
  inside[floor_65,bedroom_64]=True
  inside[window_275,home_office_246]=True
  inside[chair_101,bedroom_64]=True
  on[ceiling_272,wall_261]=True
  inside[broom_2000,bedroom_64]=True
  inside[broom_2000,dresser_100]=True
  inside[controller_2036,home_office_246]=True
  inside[faucet_29,bathroom_1]=True
  facing[powersocket_201,drawing_197]=True
  inside[wall_13,bathroom_1]=True
  inside[pillow_310,home_office_246]=True
  close[blender_2003,filing_cabinet_305]=True
  facing[tablelamp_95,drawing_110]=True
  inside[bag_2061,bedroom_64]=True
  inside[bag_2061,dresser_100]=True
  inside[drawing_110,bedroom_64]=True
  inside[wall_258,home_office_246]=True
  close[wall_175,walllamp_25]=True
  close[wall_175,floor_167]=True
  close[wall_175,floor_169]=True
  close[wall_175,floor_170]=True
  close[wall_175,wall_172]=True
  close[wall_175,wall_176]=True
  close[wall_175,ceiling_179]=True
  close[wall_175,ceiling_180]=True
  close[wall_175,ceiling_181]=True
  close[wall_175,door_183]=True
  close[wall_175,ceilinglamp_186]=True
  close[wall_175,table_189]=True
  close[wall_175,bench_190]=True
  close[wall_175,bookshelf_195]=True
  close[wall_175,mat_196]=True
  close[wall_175,drawing_198]=True
  close[wall_175,orchid_199]=True
  close[wall_175,floor_74]=True
  close[wall_175,wall_76]=True
  close[wall_175,phone_205]=True
  close[wall_175,wall_81]=True
  close[wall_175,ceiling_93]=True
  close[wall_175,cutting_board_223]=True
  close[wall_175,doorjamb_104]=True
  close[wall_175,drawing_110]=True
  close[ceiling_93,drawing_198]=True
  close[ceiling_93,doorjamb_104]=True
  close[ceiling_93,drawing_108]=True
  close[ceiling_93,phone_205]=True
  close[ceiling_93,drawing_110]=True
  close[ceiling_93,ceiling_15]=True
  close[ceiling_93,wall_12]=True
  close[ceiling_93,wall_81]=True
  close[ceiling_93,wall_175]=True
  close[ceiling_93,ceiling_180]=True
  close[ceiling_93,ceiling_88]=True
  close[ceiling_93,walllamp_25]=True
  close[ceiling_93,ceiling_92]=True
  close[ceiling_93,light_62]=True
  close[ceiling_93,towel_rack_31]=True
  on[mousepad_319,desk_282]=True
  close[ceiling_180,bookshelf_195]=True
  close[ceiling_180,drawing_198]=True
  close[ceiling_180,doorjamb_104]=True
  close[ceiling_180,wall_172]=True
  close[ceiling_180,phone_205]=True
  close[ceiling_180,drawing_110]=True
  close[ceiling_180,wall_175]=True
  close[ceiling_180,wall_81]=True
  close[ceiling_180,ceiling_179]=True
  close[ceiling_180,ceiling_181]=True
  close[ceiling_180,walllamp_25]=True
  close[ceiling_180,ceilinglamp_186]=True
  close[ceiling_180,ceiling_93]=True
  inside[check_2045,dining_room_163]=True
  close[ground_coffee_2046,filing_cabinet_305]=True
  facing[ceiling_85,drawing_109]=True
  facing[wall_257,computer_321]=True
  inside[floor_68,bedroom_64]=True
  inside[curtain_22,bathroom_1]=True
  inside[ceiling_16,bathroom_1]=True
  close[bathtub_30,towel_rack_32]=True
  close[bathtub_30,floor_5]=True
  close[bathtub_30,shelf_38]=True
  close[bathtub_30,floor_8]=True
  close[bathtub_30,wall_10]=True
  close[bathtub_30,wall_13]=True
  close[bathtub_30,curtain_22]=True
  close[bathtub_30,window_61]=True
  close[shower_35,chair_96]=True
  close[shower_35,wall_258]=True
  close[shower_35,wall_259]=True
  close[shower_35,toilet_37]=True
  close[shower_35,floor_7]=True
  close[shower_35,floor_72]=True
  close[shower_35,ceiling_264]=True
  close[shower_35,wall_11]=True
  close[shower_35,ceiling_17]=True
  close[shower_35,wall_82]=True
  close[shower_35,wall_83]=True
  close[shower_35,doorjamb_273]=True
  close[shower_35,floor_247]=True
  close[shower_35,bookshelf_280]=True
  close[shower_35,walllamp_26]=True
  close[shower_35,ceiling_91]=True
  inside[coffe_maker_236,dining_room_163]=True
  facing[ceilinglamp_187,television_202]=True
  facing[ceilinglamp_187,wall_clock_204]=True
  close[deck_of_cards_2041,dresser_100]=True
  inside[wall_77,bedroom_64]=True
  close[ceiling_178,light_200]=True
  close[ceiling_178,wall_171]=True
  close[ceiling_178,wall_172]=True
  close[ceiling_178,wall_173]=True
  close[ceiling_178,ceiling_177]=True
  close[ceiling_178,ceiling_179]=True
  close[ceiling_178,ceiling_181]=True
  close[ceiling_178,doorjamb_184]=True
  close[ceiling_178,maindoor_185]=True
  close[ceiling_178,ceilinglamp_186]=True
  close[ceiling_178,ceilinglamp_187]=True
  on[shelf_38,floor_8]=True
  close[sink_193,kitchen_counter_192]=True
  close[sink_193,faucet_194]=True
  close[sink_193,floor_164]=True
  close[sink_193,floor_165]=True
  close[sink_193,cutting_board_228]=True
  close[sink_193,toaster_231]=True
  close[sink_193,floor_166]=True
  close[sink_193,coffe_maker_236]=True
  close[sink_193,wall_173]=True
  close[sink_193,microwave_238]=True
  close[sink_193,wall_174]=True
  close[orchid_199,mat_196]=True
  close[orchid_199,floor_167]=True
  close[orchid_199,floor_168]=True
  close[orchid_199,wall_172]=True
  close[orchid_199,wall_173]=True
  close[orchid_199,wall_174]=True
  close[orchid_199,wall_175]=True
  close[orchid_199,table_189]=True
  close[orchid_199,bench_190]=True
  close[orchid_199,bench_191]=True
  close[bookshelf_280,chair_96]=True
  close[bookshelf_280,wall_258]=True
  close[bookshelf_280,wall_259]=True
  close[bookshelf_280,shower_35]=True
  close[bookshelf_280,toilet_37]=True
  close[bookshelf_280,floor_7]=True
  close[bookshelf_280,ceiling_264]=True
  close[bookshelf_280,floor_72]=True
  close[bookshelf_280,stamp_2056]=True
  close[bookshelf_280,wall_11]=True
  close[bookshelf_280,ceiling_269]=True
  close[bookshelf_280,doorjamb_273]=True
  close[bookshelf_280,wall_82]=True
  close[bookshelf_280,wall_83]=True
  close[bookshelf_280,drawing_309]=True
  close[bookshelf_280,light_316]=True
  close[bookshelf_280,floor_247]=True
  close[bookshelf_280,walllamp_26]=True
  close[bookshelf_280,floor_252]=True
  close[bookshelf_280,powersocket_317]=True
  inside[glue_2012,home_office_246]=True
  inside[wall_261,home_office_246]=True
  inside[wall_174,dining_room_163]=True
  inside[walllamp_25,bathroom_1]=True
  facing[ceiling_266,television_315]=True
  facing[ceiling_266,drawing_307]=True
  between[doorjamb_273,bedroom_64]=True
  between[doorjamb_273,home_office_246]=True
  inside[wall_9,bathroom_1]=True
  inside[food_salt_2057,bathroom_1]=True
  inside[food_salt_2057,sink_28]=True
  on[faucet_194,kitchen_counter_192]=True
  close[clothes_pants_2002,couch_279]=True
  close[comb_2017,bathroom_counter_27]=True
  inside[sink_193,kitchen_counter_192]=True
  inside[sink_193,dining_room_163]=True
  facing[mat_196,drawing_197]=True
  facing[mat_196,drawing_198]=True
  inside[oven_229,dining_room_163]=True
  inside[ceiling_270,home_office_246]=True
  close[novel_2042,desk_282]=True
  close[floor_73,floor_6]=True
  close[floor_73,door_39]=True
  close[floor_73,doorjamb_40]=True
  close[floor_73,light_105]=True
  close[floor_73,table_103]=True
  close[floor_73,floor_70]=True
  close[floor_73,floor_74]=True
  close[floor_73,floor_72]=True
  close[floor_73,wall_14]=True
  close[floor_73,wall_80]=True
  close[floor_73,wall_81]=True
  close[floor_73,light_62]=True
  close[floor_73,towel_rack_31]=True
  close[ground_coffee_1004,freezer_234]=True
  close[ceilinglamp_94,vase_115]=True
  close[ceilinglamp_94,ceiling_86]=True
  close[ceilinglamp_94,ceiling_88]=True
  close[ceilinglamp_94,ceiling_89]=True
  close[ceilinglamp_94,ceiling_90]=True
  close[ceilinglamp_94,ceiling_92]=True
  on[clothes_pants_2002,couch_279]=True
  on[pillow_2006,bench_191]=True
  inside[ceiling_177,dining_room_163]=True
  facing[floor_73,drawing_108]=True
  facing[floor_73,drawing_110]=True
  close[hanger_293,hanger_289]=True
  close[hanger_293,hanger_291]=True
  close[hanger_293,wall_260]=True
  close[hanger_293,wall_262]=True
  close[hanger_293,hanger_295]=True
  close[hanger_293,closetdrawer_296]=True
  close[hanger_293,ceiling_265]=True
  close[hanger_293,ceiling_266]=True
  close[hanger_293,closetdrawer_299]=True
  close[hanger_293,closetdrawer_301]=True
  close[hanger_293,drawing_307]=True
  close[hanger_293,dresser_284]=True
  close[hanger_293,hanger_285]=True
  close[hanger_293,hanger_287]=True
  close[closetdrawer_299,hanger_289]=True
  close[closetdrawer_299,hanger_291]=True
  close[closetdrawer_299,wall_260]=True
  close[closetdrawer_299,hanger_293]=True
  close[closetdrawer_299,hanger_295]=True
  close[closetdrawer_299,closetdrawer_296]=True
  close[closetdrawer_299,closetdrawer_301]=True
  close[closetdrawer_299,standingmirror_306]=True
  close[closetdrawer_299,floor_249]=True
  close[closetdrawer_299,dresser_284]=True
  close[closetdrawer_299,hanger_285]=True
  close[closetdrawer_299,hanger_287]=True
  facing[bookshelf_97,drawing_108]=True
  inside[closetdrawer_141,bedroom_64]=True
  inside[closetdrawer_141,dresser_100]=True
  close[broom_2049,floor_164]=True
  close[mat_21,floor_2]=True
  close[mat_21,floor_3]=True
  close[mat_21,floor_4]=True
  close[mat_21,oven_229]=True
  close[mat_21,tray_230]=True
  close[mat_21,floor_167]=True
  close[mat_21,floor_6]=True
  close[mat_21,wall_9]=True
  close[mat_21,floor_166]=True
  close[mat_21,floor_5]=True
  close[mat_21,wall_12]=True
  close[mat_21,wall_174]=True
  close[mat_21,wall_176]=True
  close[mat_21,bathroom_counter_27]=True
  close[mat_21,sink_28]=True
  close[mat_21,faucet_29]=True
  inside[microwave_238,dining_room_163]=True
  close[walllamp_26,shower_35]=True
  close[walllamp_26,wall_259]=True
  close[walllamp_26,floor_7]=True
  close[walllamp_26,ceiling_264]=True
  close[walllamp_26,floor_8]=True
  close[walllamp_26,wall_10]=True
  close[walllamp_26,wall_11]=True
  close[walllamp_26,ceiling_17]=True
  close[walllamp_26,ceiling_18]=True
  close[walllamp_26,floor_247]=True
  close[walllamp_26,bookshelf_280]=True
  inside[ceilinglamp_186,dining_room_163]=True
  on[cpuscreen_320,desk_282]=True
  close[floor_74,floor_2]=True
  close[floor_74,floor_3]=True
  close[floor_74,floor_69]=True
  close[floor_74,door_39]=True
  close[floor_74,doorjamb_104]=True
  close[floor_74,floor_73]=True
  close[floor_74,floor_170]=True
  close[floor_74,drawing_108]=True
  close[floor_74,phone_205]=True
  close[floor_74,drawing_110]=True
  close[floor_74,wall_12]=True
  close[floor_74,wall_175]=True
  close[floor_74,wall_81]=True
  close[floor_74,door_183]=True
  close[floor_74,walllamp_25]=True
  close[floor_74,light_62]=True
  close[floor_74,towel_rack_31]=True
  close[wall_80,floor_6]=True
  close[wall_80,door_39]=True
  close[wall_80,doorjamb_40]=True
  close[wall_80,light_105]=True
  close[wall_80,floor_73]=True
  close[wall_80,wall_11]=True
  close[wall_80,drawing_108]=True
  close[wall_80,wall_12]=True
  close[wall_80,wall_14]=True
  close[wall_80,ceiling_16]=True
  close[wall_80,wall_81]=True
  close[wall_80,wall_82]=True
  close[wall_80,ceiling_92]=True
  close[wall_80,light_62]=True
  close[wall_80,towel_rack_31]=True
  inside[mat_196,dining_room_163]=True
  on[bookshelf_195,floor_170]=True
  on[sheets_2058,bed_99]=True
  inside[closetdrawer_144,bedroom_64]=True
  inside[closetdrawer_144,dresser_100]=True
  close[sink_28,floor_2]=True
  close[sink_28,floor_3]=True
  close[sink_28,bathroom_cabinet_36]=True
  close[sink_28,oven_229]=True
  close[sink_28,tray_230]=True
  close[sink_28,floor_4]=True
  close[sink_28,floor_166]=True
  close[sink_28,wall_9]=True
  close[sink_28,floor_167]=True
  close[sink_28,stovefan_235]=True
  close[sink_28,wall_clock_204]=True
  close[sink_28,wall_12]=True
  close[sink_28,wall_174]=True
  close[sink_28,food_salt_2057]=True
  close[sink_28,wall_176]=True
  close[sink_28,mat_21]=True
  close[sink_28,bathroom_counter_27]=True
  close[sink_28,faucet_29]=True
  close[closetdrawer_142,wall_257]=True
  close[closetdrawer_142,hanger_130]=True
  close[closetdrawer_142,hanger_131]=True
  close[closetdrawer_142,hanger_132]=True
  close[closetdrawer_142,hanger_133]=True
  close[closetdrawer_142,hanger_134]=True
  close[closetdrawer_142,closetdrawer_141]=True
  close[closetdrawer_142,closetdrawer_143]=True
  close[closetdrawer_142,closetdrawer_144]=True
  close[closetdrawer_142,closetdrawer_145]=True
  close[closetdrawer_142,closetdrawer_146]=True
  close[closetdrawer_142,desk_282]=True
  close[closetdrawer_142,mouse_318]=True
  close[closetdrawer_142,mousepad_319]=True
  close[closetdrawer_142,cpuscreen_320]=True
  close[closetdrawer_142,computer_321]=True
  close[closetdrawer_142,keyboard_322]=True
  close[closetdrawer_142,floor_66]=True
  close[closetdrawer_142,floor_65]=True
  close[closetdrawer_142,floor_71]=True
  close[closetdrawer_142,wall_75]=True
  close[closetdrawer_142,wall_78]=True
  close[closetdrawer_142,dresser_100]=True
  close[closetdrawer_142,hanger_124]=True
  close[closetdrawer_142,floor_253]=True
  close[closetdrawer_142,hanger_126]=True
  close[closetdrawer_142,hanger_127]=True
  inside[phone_205,dining_room_163]=True
  between[door_39,bedroom_64]=True
  between[door_39,bathroom_1]=True
  on[ceiling_93,wall_81]=True
  close[hanger_132,hanger_128]=True
  close[hanger_132,hanger_129]=True
  close[hanger_132,hanger_130]=True
  close[hanger_132,hanger_131]=True
  close[hanger_132,wall_257]=True
  close[hanger_132,hanger_133]=True
  close[hanger_132,hanger_134]=True
  close[hanger_132,closetdrawer_141]=True
  close[hanger_132,closetdrawer_142]=True
  close[hanger_132,closetdrawer_143]=True
  close[hanger_132,closetdrawer_144]=True
  close[hanger_132,ceiling_270]=True
  close[hanger_132,desk_282]=True
  close[hanger_132,cpuscreen_320]=True
  close[hanger_132,keyboard_322]=True
  close[hanger_132,wall_75]=True
  close[hanger_132,wall_78]=True
  close[hanger_132,ceiling_85]=True
  close[hanger_132,ceiling_90]=True
  close[hanger_132,dresser_100]=True
  close[hanger_132,hanger_124]=True
  close[hanger_132,hanger_125]=True
  close[hanger_132,hanger_126]=True
  close[hanger_132,hanger_127]=True
  facing[doorjamb_184,drawing_197]=True
  close[ceiling_85,hanger_132]=True
  close[ceiling_85,chair_101]=True
  close[ceiling_85,hanger_134]=True
  close[ceiling_85,hanger_133]=True
  close[ceiling_85,drawing_109]=True
  close[ceiling_85,wall_78]=True
  close[ceiling_85,ceiling_86]=True
  close[ceiling_85,ceiling_90]=True
  close[ceiling_85,hanger_124]=True
  inside[curtain_112,bedroom_64]=True
  inside[curtain_112,curtain_111]=True
  facing[curtain_311,television_315]=True
  inside[milk_1003,freezer_234]=True
  inside[milk_1003,dining_room_163]=True
  inside[table_189,dining_room_163]=True
  close[curtain_311,wall_256]=True
  close[curtain_311,wall_261]=True
  close[curtain_311,ceiling_267]=True
  close[curtain_311,ceiling_272]=True
  close[curtain_311,window_275]=True
  close[curtain_311,mat_308]=True
  close[curtain_311,couch_279]=True
  close[curtain_311,curtain_312]=True
  close[curtain_311,curtain_313]=True
  close[curtain_311,floor_250]=True
  facing[bench_190,television_202]=True
  facing[bench_190,drawing_197]=True
  facing[bench_190,drawing_198]=True
  facing[curtain_313,television_315]=True
  facing[curtain_313,drawing_307]=True
  facing[floor_68,drawing_110]=True
  on[blow_dryer_2059,bathroom_counter_27]=True
  facing[ceiling_92,drawing_108]=True
  facing[ceiling_92,drawing_110]=True
  close[closetdrawer_145,cpuscreen_320]=True
  close[closetdrawer_145,computer_321]=True
  close[closetdrawer_145,keyboard_322]=True
  close[closetdrawer_145,wall_257]=True
  close[closetdrawer_145,dresser_100]=True
  close[closetdrawer_145,floor_66]=True
  close[closetdrawer_145,floor_65]=True
  close[closetdrawer_145,floor_71]=True
  close[closetdrawer_145,wall_75]=True
  close[closetdrawer_145,closetdrawer_141]=True
  close[closetdrawer_145,closetdrawer_142]=True
  close[closetdrawer_145,closetdrawer_143]=True
  close[closetdrawer_145,closetdrawer_144]=True
  close[closetdrawer_145,wall_78]=True
  close[closetdrawer_145,closetdrawer_146]=True
  close[closetdrawer_145,desk_282]=True
  close[closetdrawer_145,floor_253]=True
  close[closetdrawer_145,mouse_318]=True
  close[closetdrawer_145,mousepad_319]=True
  inside[filing_cabinet_305,home_office_246]=True
  close[ceiling_87,bookshelf_97]=True
  close[ceiling_87,hanger_102]=True
  close[ceiling_87,curtain_111]=True
  close[ceiling_87,curtain_112]=True
  close[ceiling_87,wall_79]=True
  close[ceiling_87,ceiling_86]=True
  close[ceiling_87,ceiling_88]=True
  inside[wall_172,dining_room_163]=True
  on[toaster_231,kitchen_counter_192]=True
  close[ceiling_92,doorjamb_40]=True
  close[ceiling_92,light_105]=True
  close[ceiling_92,drawing_108]=True
  close[ceiling_92,wall_14]=True
  close[ceiling_92,wall_80]=True
  close[ceiling_92,ceiling_16]=True
  close[ceiling_92,wall_81]=True
  close[ceiling_92,ceilinglamp_94]=True
  close[ceiling_92,ceiling_89]=True
  close[ceiling_92,ceiling_91]=True
  close[ceiling_92,ceiling_93]=True
  close[ceiling_92,light_62]=True
  close[ceiling_92,towel_rack_31]=True
  close[floor_170,bookshelf_195]=True
  close[floor_170,floor_167]=True
  close[floor_170,doorjamb_104]=True
  close[floor_170,floor_169]=True
  close[floor_170,floor_74]=True
  close[floor_170,wall_172]=True
  close[floor_170,phone_205]=True
  close[floor_170,drawing_110]=True
  close[floor_170,wall_175]=True
  close[floor_170,wall_81]=True
  close[floor_170,door_183]=True
  close[floor_170,walllamp_25]=True
  close[floor_170,table_189]=True
  close[floor_170,bench_190]=True
  close[floor_170,cutting_board_223]=True
  close[maindoor_185,floor_168]=True
  close[maindoor_185,powersocket_201]=True
  close[maindoor_185,light_200]=True
  close[maindoor_185,wall_171]=True
  close[maindoor_185,wall_172]=True
  close[maindoor_185,wall_173]=True
  close[maindoor_185,ceiling_178]=True
  close[maindoor_185,doorjamb_184]=True
  on[photoframe_219,tvstand_188]=True
  inside[tablelamp_95,bedroom_64]=True
  inside[clothes_pants_2040,bedroom_64]=True
  inside[clothes_pants_2040,dresser_100]=True
  on[door_183,floor_74]=True
  on[mouthwash_2027,bathroom_counter_27]=True
  close[floor_254,wall_257]=True
  close[floor_254,wall_261]=True
  close[floor_254,wall_263]=True
  close[floor_254,piano_bench_2047]=True
  close[floor_254,floor_251]=True
  close[floor_254,television_315]=True
  close[floor_254,doorjamb_274]=True
  close[floor_254,mat_308]=True
  close[floor_254,piano_bench_2005]=True
  close[floor_254,walllamp_278]=True
  close[floor_254,couch_279]=True
  close[floor_254,table_281]=True
  close[floor_254,chair_283]=True
  close[floor_254,floor_253]=True
  close[floor_254,floor_255]=True
  inside[fork_2004,home_office_246]=True
  inside[toy_314,home_office_246]=True
  facing[wall_263,computer_321]=True
  facing[wall_263,television_315]=True
  close[broom_2000,dresser_100]=True
  close[food_food_2009,table_103]=True
  close[juice_1006,freezer_234]=True
  close[closetdrawer_141,hanger_128]=True
  close[closetdrawer_141,hanger_129]=True
  close[closetdrawer_141,hanger_130]=True
  close[closetdrawer_141,hanger_131]=True
  close[closetdrawer_141,hanger_132]=True
  close[closetdrawer_141,hanger_133]=True
  close[closetdrawer_141,hanger_134]=True
  close[closetdrawer_141,wall_257]=True
  close[closetdrawer_141,closetdrawer_142]=True
  close[closetdrawer_141,closetdrawer_143]=True
  close[closetdrawer_141,closetdrawer_144]=True
  close[closetdrawer_141,closetdrawer_145]=True
  close[closetdrawer_141,closetdrawer_146]=True
  close[closetdrawer_141,desk_282]=True
  close[closetdrawer_141,mouse_318]=True
  close[closetdrawer_141,mousepad_319]=True
  close[closetdrawer_141,cpuscreen_320]=True
  close[closetdrawer_141,computer_321]=True
  close[closetdrawer_141,keyboard_322]=True
  close[closetdrawer_141,floor_66]=True
  close[closetdrawer_141,floor_65]=True
  close[closetdrawer_141,floor_71]=True
  close[closetdrawer_141,wall_75]=True
  close[closetdrawer_141,wall_78]=True
  close[closetdrawer_141,dresser_100]=True
  close[closetdrawer_141,floor_253]=True
  close[closetdrawer_141,hanger_124]=True
  close[closetdrawer_141,hanger_125]=True
  close[closetdrawer_141,hanger_126]=True
  close[closetdrawer_141,hanger_127]=True
  facing[window_275,television_315]=True
  close[closetdrawer_146,wall_257]=True
  close[closetdrawer_146,wall_258]=True
  close[closetdrawer_146,closetdrawer_141]=True
  close[closetdrawer_146,closetdrawer_142]=True
  close[closetdrawer_146,closetdrawer_143]=True
  close[closetdrawer_146,closetdrawer_144]=True
  close[closetdrawer_146,closetdrawer_145]=True
  close[closetdrawer_146,desk_282]=True
  close[closetdrawer_146,light_316]=True
  close[closetdrawer_146,powersocket_317]=True
  close[closetdrawer_146,mouse_318]=True
  close[closetdrawer_146,mousepad_319]=True
  close[closetdrawer_146,cpuscreen_320]=True
  close[closetdrawer_146,computer_321]=True
  close[closetdrawer_146,keyboard_322]=True
  close[closetdrawer_146,floor_71]=True
  close[closetdrawer_146,floor_72]=True
  close[closetdrawer_146,wall_75]=True
  close[closetdrawer_146,wall_83]=True
  close[closetdrawer_146,dresser_100]=True
  close[closetdrawer_146,floor_252]=True
  close[closetdrawer_146,floor_253]=True
  inside[ceiling_88,bedroom_64]=True
  close[clothes_pants_2040,dresser_100]=True
  inside[hanger_124,bedroom_64]=True
  inside[hanger_124,dresser_100]=True
  inside[floor_165,dining_room_163]=True
  facing[closetdrawer_299,television_315]=True
  inside[video_game_controller_2039,dining_room_163]=True
  inside[ceiling_272,home_office_246]=True
  close[kitchen_counter_192,food_carrot_2016]=True
  close[kitchen_counter_192,sink_193]=True
  close[kitchen_counter_192,faucet_194]=True
  close[kitchen_counter_192,floor_164]=True
  close[kitchen_counter_192,floor_165]=True
  close[kitchen_counter_192,cutting_board_228]=True
  close[kitchen_counter_192,toaster_231]=True
  close[kitchen_counter_192,floor_166]=True
  close[kitchen_counter_192,tray_230]=True
  close[kitchen_counter_192,freezer_234]=True
  close[kitchen_counter_192,oven_229]=True
  close[kitchen_counter_192,coffe_maker_236]=True
  close[kitchen_counter_192,wall_173]=True
  close[kitchen_counter_192,microwave_238]=True
  close[kitchen_counter_192,wall_174]=True
  close[kitchen_counter_192,food_rice_2038]=True
  close[kitchen_counter_192,cup_2008]=True
  close[kitchen_counter_192,towel_2011]=True
  facing[floor_166,wall_clock_204]=True
  close[hanger_291,hanger_289]=True
  close[hanger_291,wall_260]=True
  close[hanger_291,hanger_293]=True
  close[hanger_291,wall_262]=True
  close[hanger_291,hanger_295]=True
  close[hanger_291,closetdrawer_296]=True
  close[hanger_291,ceiling_265]=True
  close[hanger_291,ceiling_266]=True
  close[hanger_291,closetdrawer_299]=True
  close[hanger_291,closetdrawer_301]=True
  close[hanger_291,drawing_307]=True
  close[hanger_291,dresser_284]=True
  close[hanger_291,hanger_285]=True
  close[hanger_291,hanger_287]=True
  inside[floor_72,bedroom_64]=True
  close[closetdrawer_296,hanger_289]=True
  close[closetdrawer_296,hanger_291]=True
  close[closetdrawer_296,wall_260]=True
  close[closetdrawer_296,hanger_293]=True
  close[closetdrawer_296,wall_262]=True
  close[closetdrawer_296,hanger_295]=True
  close[closetdrawer_296,closetdrawer_299]=True
  close[closetdrawer_296,closetdrawer_301]=True
  close[closetdrawer_296,standingmirror_306]=True
  close[closetdrawer_296,drawing_307]=True
  close[closetdrawer_296,floor_248]=True
  close[closetdrawer_296,floor_249]=True
  close[closetdrawer_296,dresser_284]=True
  close[closetdrawer_296,hanger_285]=True
  close[closetdrawer_296,hanger_287]=True
  inside[laundry_detergent_2023,filing_cabinet_305]=True
  inside[laundry_detergent_2023,home_office_246]=True
  close[floor_249,wall_260]=True
  close[floor_249,closetdrawer_296]=True
  close[floor_249,closetdrawer_299]=True
  close[floor_249,closetdrawer_301]=True
  close[floor_249,standingmirror_306]=True
  close[floor_249,floor_248]=True
  close[floor_249,floor_250]=True
  close[floor_249,dresser_284]=True
  inside[bathroom_cabinet_36,bathroom_1]=True
  facing[wall_80,drawing_110]=True
  inside[table_281,home_office_246]=True
  inside[mat_107,bedroom_64]=True
  inside[powersocket_317,home_office_246]=True
  close[floor_72,wall_258]=True
  close[floor_72,floor_7]=True
  close[floor_72,wall_11]=True
  close[floor_72,closetdrawer_143]=True
  close[floor_72,closetdrawer_144]=True
  close[floor_72,doorjamb_273]=True
  close[floor_72,closetdrawer_146]=True
  close[floor_72,bookshelf_280]=True
  close[floor_72,desk_282]=True
  close[floor_72,shower_35]=True
  close[floor_72,toilet_37]=True
  close[floor_72,door_39]=True
  close[floor_72,light_316]=True
  close[floor_72,powersocket_317]=True
  close[floor_72,mouse_318]=True
  close[floor_72,mousepad_319]=True
  close[floor_72,computer_321]=True
  close[floor_72,floor_71]=True
  close[floor_72,floor_73]=True
  close[floor_72,wall_82]=True
  close[floor_72,wall_83]=True
  close[floor_72,chair_96]=True
  close[floor_72,light_105]=True
  close[floor_72,floor_252]=True
  close[ceiling_267,wall_256]=True
  close[ceiling_267,wall_260]=True
  close[ceiling_267,wall_261]=True
  close[ceiling_267,ceiling_266]=True
  close[ceiling_267,ceiling_268]=True
  close[ceiling_267,ceiling_272]=True
  close[ceiling_267,standingmirror_306]=True
  close[ceiling_267,window_275]=True
  close[ceiling_267,ceilinglamp_276]=True
  close[ceiling_267,curtain_311]=True
  close[ceiling_267,curtain_312]=True
  close[ceiling_267,curtain_313]=True
  inside[floor_71,bedroom_64]=True
  inside[food_carrot_2016,dining_room_163]=True
  inside[ceiling_265,home_office_246]=True
  inside[ceiling_91,bedroom_64]=True
  inside[hanger_132,bedroom_64]=True
  inside[hanger_132,dresser_100]=True
  close[phone_205,floor_2]=True
  close[phone_205,floor_3]=True
  close[phone_205,bathroom_cabinet_36]=True
  close[phone_205,floor_167]=True
  close[phone_205,doorjamb_104]=True
  close[phone_205,floor_170]=True
  close[phone_205,floor_74]=True
  close[phone_205,wall_clock_204]=True
  close[phone_205,wall_12]=True
  close[phone_205,drawing_108]=True
  close[phone_205,ceiling_15]=True
  close[phone_205,wall_176]=True
  close[phone_205,wall_175]=True
  close[phone_205,wall_81]=True
  close[phone_205,ceiling_180]=True
  close[phone_205,ceiling_181]=True
  close[phone_205,door_183]=True
  close[phone_205,walllamp_25]=True
  close[phone_205,bathroom_counter_27]=True
  close[phone_205,ceiling_93]=True
  facing[maindoor_185,drawing_197]=True
  inside[check_2026,filing_cabinet_305]=True
  inside[check_2026,home_office_246]=True
  close[coffe_maker_236,kitchen_counter_192]=True
  close[coffe_maker_236,sink_193]=True
  close[coffe_maker_236,faucet_194]=True
  close[coffe_maker_236,cutting_board_228]=True
  close[coffe_maker_236,floor_165]=True
  close[coffe_maker_236,floor_164]=True
  close[coffe_maker_236,toaster_231]=True
  close[coffe_maker_236,floor_166]=True
  close[coffe_maker_236,freezer_234]=True
  close[coffe_maker_236,wall_173]=True
  close[coffe_maker_236,microwave_238]=True
  close[coffe_maker_236,wall_174]=True
  close[coffe_maker_236,ceiling_177]=True
  close[coffe_maker_236,ceiling_182]=True
  close[floor_251,mat_308]=True
  close[floor_251,couch_279]=True
  close[floor_251,floor_248]=True
  close[floor_251,table_281]=True
  close[floor_251,floor_250]=True
  close[floor_251,television_315]=True
  close[floor_251,floor_252]=True
  close[floor_251,floor_254]=True
  close[blender_2048,cupboard_1000]=True
  close[ceiling_20,towel_rack_33]=True
  close[ceiling_20,wallshelf_34]=True
  close[ceiling_20,bathroom_cabinet_36]=True
  close[ceiling_20,wall_9]=True
  close[ceiling_20,stovefan_235]=True
  close[ceiling_20,wall_clock_204]=True
  close[ceiling_20,wall_12]=True
  close[ceiling_20,wall_174]=True
  close[ceiling_20,ceiling_15]=True
  close[ceiling_20,ceiling_19]=True
  close[ceiling_20,ceiling_182]=True
  close[ceiling_20,ceilinglamp_23]=True
  close[ceiling_20,walllamp_24]=True
  close[ceiling_20,curtain_22]=True
  close[ceiling_20,faucet_29]=True
  facing[wall_79,drawing_110]=True
  close[shaving_cream_2007,bathroom_counter_27]=True
  inside[floor_3,bathroom_1]=True
  inside[check_2051,filing_cabinet_305]=True
  inside[check_2051,home_office_246]=True
  close[glue_2012,desk_282]=True
  inside[cpuscreen_320,home_office_246]=True
  facing[table_103,drawing_108]=True
  facing[table_103,drawing_109]=True
  facing[table_103,drawing_110]=True
  inside[dresser_100,bedroom_64]=True
  facing[vase_115,drawing_108]=True
  facing[vase_115,drawing_109]=True
  facing[vase_115,drawing_110]=True
  close[wall_257,hanger_128]=True
  close[wall_257,hanger_129]=True
  close[wall_257,hanger_130]=True
  close[wall_257,hanger_131]=True
  close[wall_257,hanger_132]=True
  close[wall_257,hanger_133]=True
  close[wall_257,hanger_134]=True
  close[wall_257,wall_258]=True
  close[wall_257,wall_263]=True
  close[wall_257,closetdrawer_141]=True
  close[wall_257,ceiling_270]=True
  close[wall_257,closetdrawer_143]=True
  close[wall_257,closetdrawer_142]=True
  close[wall_257,closetdrawer_144]=True
  close[wall_257,closetdrawer_145]=True
  close[wall_257,closetdrawer_146]=True
  close[wall_257,doorjamb_274]=True
  close[wall_257,ceiling_269]=True
  close[wall_257,walllamp_278]=True
  close[wall_257,ceiling_271]=True
  close[wall_257,doorjamb_273]=True
  close[wall_257,desk_282]=True
  close[wall_257,chair_283]=True
  close[wall_257,light_316]=True
  close[wall_257,powersocket_317]=True
  close[wall_257,mouse_318]=True
  close[wall_257,mousepad_319]=True
  close[wall_257,cpuscreen_320]=True
  close[wall_257,computer_321]=True
  close[wall_257,keyboard_322]=True
  close[wall_257,floor_71]=True
  close[wall_257,wall_75]=True
  close[wall_257,wall_83]=True
  close[wall_257,ceiling_90]=True
  close[wall_257,dresser_100]=True
  close[wall_257,floor_252]=True
  close[wall_257,hanger_125]=True
  close[wall_257,floor_254]=True
  close[wall_257,hanger_124]=True
  close[wall_257,floor_253]=True
  close[wall_257,hanger_126]=True
  close[wall_257,hanger_127]=True
  close[walllamp_278,wall_257]=True
  close[walllamp_278,wall_263]=True
  close[walllamp_278,ceiling_270]=True
  close[walllamp_278,ceiling_271]=True
  close[walllamp_278,doorjamb_274]=True
  close[walllamp_278,desk_282]=True
  close[walllamp_278,chair_283]=True
  close[walllamp_278,floor_253]=True
  close[walllamp_278,floor_254]=True
  inside[dresser_284,home_office_246]=True
  inside[fork_2035,cupboard_1000]=True
  inside[fork_2035,dining_room_163]=True
  facing[floor_69,drawing_108]=True
  facing[floor_69,drawing_110]=True
  close[desk_282,hanger_128]=True
  close[desk_282,wall_257]=True
  close[desk_282,hanger_130]=True
  close[desk_282,hanger_131]=True
  close[desk_282,hanger_132]=True
  close[desk_282,hanger_133]=True
  close[desk_282,hanger_134]=True
  close[desk_282,hanger_129]=True
  close[desk_282,wall_258]=True
  close[desk_282,closetdrawer_141]=True
  close[desk_282,closetdrawer_142]=True
  close[desk_282,closetdrawer_143]=True
  close[desk_282,closetdrawer_144]=True
  close[desk_282,closetdrawer_145]=True
  close[desk_282,closetdrawer_146]=True
  close[desk_282,doorjamb_273]=True
  close[desk_282,walllamp_278]=True
  close[desk_282,chair_283]=True
  close[desk_282,light_316]=True
  close[desk_282,powersocket_317]=True
  close[desk_282,mouse_318]=True
  close[desk_282,mousepad_319]=True
  close[desk_282,cpuscreen_320]=True
  close[desk_282,computer_321]=True
  close[desk_282,keyboard_322]=True
  close[desk_282,floor_71]=True
  close[desk_282,floor_72]=True
  close[desk_282,wall_75]=True
  close[desk_282,wall_83]=True
  close[desk_282,fork_2004]=True
  close[desk_282,glue_2012]=True
  close[desk_282,dresser_100]=True
  close[desk_282,floor_252]=True
  close[desk_282,hanger_125]=True
  close[desk_282,novel_2042]=True
  close[desk_282,hanger_124]=True
  close[desk_282,floor_253]=True
  close[desk_282,hanger_126]=True
  close[desk_282,hanger_127]=True
  on[mat_196,table_189]=True
  inside[window_84,bedroom_64]=True
  facing[ceiling_93,drawing_108]=True
  facing[ceiling_93,drawing_110]=True
  close[filing_cabinet_305,wall_259]=True
  close[filing_cabinet_305,check_2051]=True
  close[filing_cabinet_305,wall_262]=True
  close[filing_cabinet_305,laundry_detergent_2023]=True
  close[filing_cabinet_305,check_2026]=True
  close[filing_cabinet_305,check_2060]=True
  close[filing_cabinet_305,needle_2030]=True
  close[filing_cabinet_305,sheets_2062]=True
  close[filing_cabinet_305,drawing_307]=True
  close[filing_cabinet_305,blender_2003]=True
  close[filing_cabinet_305,walllamp_277]=True
  close[filing_cabinet_305,drawing_309]=True
  close[filing_cabinet_305,floor_247]=True
  close[filing_cabinet_305,floor_248]=True
  close[filing_cabinet_305,centerpiece_2037]=True
  close[filing_cabinet_305,toy_314]=True
  close[filing_cabinet_305,ground_coffee_2046]=True
  close[filing_cabinet_305,drawing_2014]=True
  inside[food_food_2019,dining_room_163]=True
  inside[food_food_2019,oven_229]=True
  inside[wall_12,bathroom_1]=True
  inside[check_2060,filing_cabinet_305]=True
  inside[check_2060,home_office_246]=True
  inside[towel_rack_32,bathroom_1]=True
  on[mouse_318,desk_282]=True
  on[mouse_318,mousepad_319]=True
  close[door_39,floor_2]=True
  close[door_39,floor_3]=True
  close[door_39,floor_6]=True
  close[door_39,floor_7]=True
  close[door_39,doorjamb_40]=True
  close[door_39,light_105]=True
  close[door_39,floor_73]=True
  close[door_39,floor_74]=True
  close[door_39,drawing_108]=True
  close[door_39,floor_72]=True
  close[door_39,wall_14]=True
  close[door_39,wall_11]=True
  close[door_39,wall_80]=True
  close[door_39,wall_81]=True
  close[door_39,wall_82]=True
  close[door_39,wall_12]=True
  close[door_39,light_62]=True
  on[ceiling_177,wall_173]=True
  inside[floor_252,home_office_246]=True
  inside[hanger_293,dresser_284]=True
  inside[hanger_293,home_office_246]=True
  on[ceiling_266,wall_260]=True
  facing[wall_14,drawing_110]=True
  on[ceiling_270,wall_257]=True
  facing[wall_171,drawing_197]=True
  close[wall_79,bookshelf_97]=True
  close[wall_79,nightstand_98]=True
  close[wall_79,bed_99]=True
  close[wall_79,floor_68]=True
  close[wall_79,floor_69]=True
  close[wall_79,hanger_102]=True
  close[wall_79,floor_67]=True
  close[wall_79,mat_107]=True
  close[wall_79,wall_76]=True
  close[wall_79,wall_77]=True
  close[wall_79,curtain_111]=True
  close[wall_79,curtain_112]=True
  close[wall_79,pillow_113]=True
  close[wall_79,pillow_114]=True
  close[wall_79,vase_115]=True
  close[wall_79,window_84]=True
  close[wall_79,ceiling_86]=True
  close[wall_79,ceiling_87]=True
  close[wall_79,ceiling_88]=True
  close[wall_79,tablelamp_95]=True
  close[window_84,nightstand_98]=True
  close[window_84,bed_99]=True
  close[window_84,floor_67]=True
  close[window_84,mat_107]=True
  close[window_84,wall_77]=True
  close[window_84,wall_78]=True
  close[window_84,curtain_111]=True
  close[window_84,curtain_112]=True
  close[window_84,pillow_113]=True
  close[window_84,pillow_114]=True
  close[window_84,wall_79]=True
  close[window_84,ceiling_86]=True
  close[window_84,tablelamp_95]=True
  on[closetdrawer_141,closetdrawer_142]=True
  inside[light_200,dining_room_163]=True
  inside[floor_67,bedroom_64]=True
  inside[walllamp_277,home_office_246]=True
  inside[clothes_pants_2002,home_office_246]=True
  inside[towel_rack_31,bathroom_1]=True
  close[computer_321,wall_257]=True
  close[computer_321,wall_258]=True
  close[computer_321,closetdrawer_141]=True
  close[computer_321,closetdrawer_142]=True
  close[computer_321,closetdrawer_143]=True
  close[computer_321,closetdrawer_144]=True
  close[computer_321,closetdrawer_145]=True
  close[computer_321,closetdrawer_146]=True
  close[computer_321,desk_282]=True
  close[computer_321,chair_283]=True
  close[computer_321,light_316]=True
  close[computer_321,powersocket_317]=True
  close[computer_321,mouse_318]=True
  close[computer_321,mousepad_319]=True
  close[computer_321,cpuscreen_320]=True
  close[computer_321,keyboard_322]=True
  close[computer_321,floor_71]=True
  close[computer_321,floor_72]=True
  close[computer_321,wall_75]=True
  close[computer_321,wall_83]=True
  close[computer_321,dresser_100]=True
  close[computer_321,floor_252]=True
  close[computer_321,floor_253]=True
  facing[doorjamb_274,computer_321]=True
  facing[doorjamb_274,television_315]=True
  on[video_game_controller_2039,table_189]=True
  inside[stovefan_235,dining_room_163]=True
  inside[ceiling_15,bathroom_1]=True
  inside[closetdrawer_296,dresser_284]=True
  inside[closetdrawer_296,home_office_246]=True
  inside[band_aids_2063,bedroom_64]=True
  inside[band_aids_2063,dresser_100]=True
  facing[ceiling_180,drawing_108]=True
  facing[ceiling_180,drawing_197]=True
  facing[ceiling_180,drawing_198]=True
  close[hanger_133,hanger_128]=True
  close[hanger_133,hanger_129]=True
  close[hanger_133,hanger_130]=True
  close[hanger_133,hanger_131]=True
  close[hanger_133,hanger_132]=True
  close[hanger_133,wall_257]=True
  close[hanger_133,hanger_134]=True
  close[hanger_133,closetdrawer_141]=True
  close[hanger_133,closetdrawer_142]=True
  close[hanger_133,closetdrawer_143]=True
  close[hanger_133,closetdrawer_144]=True
  close[hanger_133,ceiling_270]=True
  close[hanger_133,desk_282]=True
  close[hanger_133,cpuscreen_320]=True
  close[hanger_133,keyboard_322]=True
  close[hanger_133,wall_75]=True
  close[hanger_133,wall_78]=True
  close[hanger_133,ceiling_85]=True
  close[hanger_133,ceiling_90]=True
  close[hanger_133,dresser_100]=True
  close[hanger_133,hanger_124]=True
  close[hanger_133,hanger_125]=True
  close[hanger_133,hanger_126]=True
  close[hanger_133,hanger_127]=True
  close[closetdrawer_144,hanger_128]=True
  close[closetdrawer_144,hanger_129]=True
  close[closetdrawer_144,hanger_130]=True
  close[closetdrawer_144,hanger_131]=True
  close[closetdrawer_144,hanger_132]=True
  close[closetdrawer_144,hanger_133]=True
  close[closetdrawer_144,hanger_134]=True
  close[closetdrawer_144,wall_257]=True
  close[closetdrawer_144,wall_258]=True
  close[closetdrawer_144,closetdrawer_141]=True
  close[closetdrawer_144,closetdrawer_142]=True
  close[closetdrawer_144,closetdrawer_143]=True
  close[closetdrawer_144,closetdrawer_145]=True
  close[closetdrawer_144,closetdrawer_146]=True
  close[closetdrawer_144,desk_282]=True
  close[closetdrawer_144,light_316]=True
  close[closetdrawer_144,powersocket_317]=True
  close[closetdrawer_144,mouse_318]=True
  close[closetdrawer_144,mousepad_319]=True
  close[closetdrawer_144,cpuscreen_320]=True
  close[closetdrawer_144,computer_321]=True
  close[closetdrawer_144,keyboard_322]=True
  close[closetdrawer_144,floor_71]=True
  close[closetdrawer_144,floor_72]=True
  close[closetdrawer_144,wall_75]=True
  close[closetdrawer_144,wall_83]=True
  close[closetdrawer_144,dresser_100]=True
  close[closetdrawer_144,floor_252]=True
  close[closetdrawer_144,floor_253]=True
  close[closetdrawer_144,hanger_124]=True
  close[closetdrawer_144,hanger_125]=True
  close[closetdrawer_144,hanger_126]=True
  close[closetdrawer_144,hanger_127]=True
  inside[photoframe_219,dining_room_163]=True
  inside[wall_260,home_office_246]=True
  facing[wall_clock_204,drawing_198]=True
  close[wall_82,chair_96]=True
  close[wall_82,wall_258]=True
  close[wall_82,shower_35]=True
  close[wall_82,wall_259]=True
  close[wall_82,toilet_37]=True
  close[wall_82,floor_7]=True
  close[wall_82,floor_72]=True
  close[wall_82,light_105]=True
  close[wall_82,doorjamb_40]=True
  close[wall_82,wall_11]=True
  close[wall_82,door_39]=True
  close[wall_82,wall_14]=True
  close[wall_82,wall_80]=True
  close[wall_82,doorjamb_273]=True
  close[wall_82,ceiling_17]=True
  close[wall_82,wall_83]=True
  close[wall_82,bookshelf_280]=True
  close[wall_82,ceiling_91]=True
  close[bookshelf_97,floor_68]=True
  close[bookshelf_97,floor_69]=True
  close[bookshelf_97,hanger_102]=True
  close[bookshelf_97,wall_76]=True
  close[bookshelf_97,form_2029]=True
  close[bookshelf_97,drawing_110]=True
  close[bookshelf_97,wall_79]=True
  close[bookshelf_97,ceiling_87]=True
  close[bookshelf_97,ceiling_88]=True
  close[doorjamb_184,light_200]=True
  close[doorjamb_184,powersocket_201]=True
  close[doorjamb_184,floor_168]=True
  close[doorjamb_184,wall_171]=True
  close[doorjamb_184,wall_172]=True
  close[doorjamb_184,wall_173]=True
  close[doorjamb_184,ceiling_178]=True
  close[doorjamb_184,maindoor_185]=True
  inside[door_183,dining_room_163]=True
  facing[wall_81,drawing_108]=True
  facing[wall_81,drawing_110]=True
  close[powersocket_317,chair_96]=True
  close[powersocket_317,computer_321]=True
  close[powersocket_317,wall_258]=True
  close[powersocket_317,wall_257]=True
  close[powersocket_317,dresser_100]=True
  close[powersocket_317,floor_71]=True
  close[powersocket_317,floor_72]=True
  close[powersocket_317,wall_75]=True
  close[powersocket_317,closetdrawer_143]=True
  close[powersocket_317,closetdrawer_144]=True
  close[powersocket_317,doorjamb_273]=True
  close[powersocket_317,closetdrawer_146]=True
  close[powersocket_317,wall_83]=True
  close[powersocket_317,floor_252]=True
  close[powersocket_317,bookshelf_280]=True
  close[powersocket_317,desk_282]=True
  close[powersocket_317,light_316]=True
  close[powersocket_317,floor_253]=True
  close[powersocket_317,mouse_318]=True
  close[powersocket_317,mousepad_319]=True
  on[tablelamp_95,nightstand_98]=True
  inside[floor_8,bathroom_1]=True
  inside[stamp_2056,home_office_246]=True
  on[video_game_controller_2028,table_103]=True
  on[food_carrot_2016,kitchen_counter_192]=True
  inside[ceiling_18,bathroom_1]=True
  inside[cutting_board_228,dining_room_163]=True
  inside[floor_248,home_office_246]=True
  inside[wall_176,dining_room_163]=True
  close[bowl_1001,cupboard_1000]=True
  close[wall_259,wall_258]=True
  close[wall_259,wall_262]=True
  close[wall_259,floor_7]=True
  close[wall_259,ceiling_264]=True
  close[wall_259,ceiling_265]=True
  close[wall_259,wall_11]=True
  close[wall_259,ceiling_269]=True
  close[wall_259,doorjamb_273]=True
  close[wall_259,ceiling_17]=True
  close[wall_259,walllamp_277]=True
  close[wall_259,bookshelf_280]=True
  close[wall_259,walllamp_26]=True
  close[wall_259,shower_35]=True
  close[wall_259,toilet_37]=True
  close[wall_259,filing_cabinet_305]=True
  close[wall_259,drawing_309]=True
  close[wall_259,toy_314]=True
  close[wall_259,wall_82]=True
  close[wall_259,wall_83]=True
  close[wall_259,chair_96]=True
  close[wall_259,floor_247]=True
  close[wall_259,floor_248]=True
  close[wall_259,floor_252]=True
  close[drawing_197,bookshelf_195]=True
  close[drawing_197,television_202]=True
  close[drawing_197,wall_172]=True
  close[drawing_197,ceiling_179]=True
  close[drawing_197,photoframe_219]=True
  close[drawing_197,tvstand_188]=True
  facing[ceiling_90,drawing_109]=True
  inside[bathroom_counter_27,bathroom_1]=True
  close[cutting_board_228,kitchen_counter_192]=True
  close[cutting_board_228,sink_193]=True
  close[cutting_board_228,faucet_194]=True
  close[cutting_board_228,oven_229]=True
  close[cutting_board_228,floor_166]=True
  close[cutting_board_228,freezer_234]=True
  close[cutting_board_228,coffe_maker_236]=True
  close[cutting_board_228,wall_173]=True
  close[cutting_board_228,wall_174]=True
  close[cutting_board_228,microwave_238]=True
  close[cutting_board_228,ceiling_177]=True
  close[cutting_board_228,ceiling_182]=True
  facing[pillow_114,drawing_109]=True
  close[floor_248,wall_259]=True
  close[floor_248,wall_260]=True
  close[floor_248,wall_262]=True
  close[floor_248,table_281]=True
  close[floor_248,closetdrawer_296]=True
  close[floor_248,closetdrawer_301]=True
  close[floor_248,filing_cabinet_305]=True
  close[floor_248,television_315]=True
  close[floor_248,floor_247]=True
  close[floor_248,floor_249]=True
  close[floor_248,toy_314]=True
  close[floor_248,floor_251]=True
  inside[floor_247,home_office_246]=True
  on[bathroom_cabinet_36,wall_12]=True
  facing[floor_168,drawing_197]=True
  facing[floor_168,drawing_198]=True
  inside[bookshelf_195,dining_room_163]=True
  close[purse_2022,couch_279]=True
  close[mouthwash_2027,bathroom_counter_27]=True
  inside[toaster_231,dining_room_163]=True
  facing[kitchen_counter_192,wall_clock_204]=True
  facing[hanger_295,television_315]=True
  close[piano_bench_2047,floor_254]=True
  close[ceiling_270,hanger_128]=True
  close[ceiling_270,wall_257]=True
  close[ceiling_270,hanger_130]=True
  close[ceiling_270,hanger_131]=True
  close[ceiling_270,hanger_132]=True
  close[ceiling_270,hanger_133]=True
  close[ceiling_270,hanger_134]=True
  close[ceiling_270,hanger_129]=True
  close[ceiling_270,ceiling_269]=True
  close[ceiling_270,ceiling_271]=True
  close[ceiling_270,walllamp_278]=True
  close[ceiling_270,chair_283]=True
  close[ceiling_270,light_316]=True
  close[ceiling_270,cpuscreen_320]=True
  close[ceiling_270,wall_75]=True
  close[ceiling_270,ceiling_90]=True
  close[ceiling_270,dresser_100]=True
  close[ceiling_270,hanger_124]=True
  close[ceiling_270,hanger_125]=True
  close[ceiling_270,hanger_126]=True
  close[ceiling_270,hanger_127]=True
  close[food_oatmeal_1002,cupboard_1000]=True
  inside[ceiling_179,dining_room_163]=True
  on[ceiling_17,wall_11]=True
  close[wall_clock_204,bathroom_cabinet_36]=True
  close[wall_clock_204,wall_9]=True
  close[wall_clock_204,stovefan_235]=True
  close[wall_clock_204,wall_12]=True
  close[wall_clock_204,phone_205]=True
  close[wall_clock_204,wall_174]=True
  close[wall_clock_204,ceiling_15]=True
  close[wall_clock_204,wall_176]=True
  close[wall_clock_204,ceiling_20]=True
  close[wall_clock_204,ceiling_181]=True
  close[wall_clock_204,ceiling_182]=True
  close[wall_clock_204,walllamp_25]=True
  close[wall_clock_204,bathroom_counter_27]=True
  close[wall_clock_204,sink_28]=True
  close[wall_clock_204,faucet_29]=True
  close[mouse_318,hanger_128]=True
  close[mouse_318,wall_257]=True
  close[mouse_318,hanger_129]=True
  close[mouse_318,hanger_130]=True
  close[mouse_318,hanger_131]=True
  close[mouse_318,wall_258]=True
  close[mouse_318,closetdrawer_141]=True
  close[mouse_318,closetdrawer_142]=True
  close[mouse_318,closetdrawer_143]=True
  close[mouse_318,closetdrawer_144]=True
  close[mouse_318,doorjamb_273]=True
  close[mouse_318,closetdrawer_146]=True
  close[mouse_318,closetdrawer_145]=True
  close[mouse_318,desk_282]=True
  close[mouse_318,chair_283]=True
  close[mouse_318,light_316]=True
  close[mouse_318,powersocket_317]=True
  close[mouse_318,mousepad_319]=True
  close[mouse_318,cpuscreen_320]=True
  close[mouse_318,computer_321]=True
  close[mouse_318,keyboard_322]=True
  close[mouse_318,floor_71]=True
  close[mouse_318,floor_72]=True
  close[mouse_318,wall_75]=True
  close[mouse_318,wall_83]=True
  close[mouse_318,dresser_100]=True
  close[mouse_318,floor_253]=True
  close[mouse_318,floor_252]=True
  close[mouse_318,hanger_125]=True
  close[mouse_318,hanger_126]=True
  close[mouse_318,hanger_127]=True
  facing[drawing_198,drawing_108]=True
  inside[closetdrawer_143,bedroom_64]=True
  inside[closetdrawer_143,dresser_100]=True
  close[floor_6,floor_2]=True
  close[floor_6,floor_3]=True
  close[floor_6,floor_5]=True
  close[floor_6,door_39]=True
  close[floor_6,doorjamb_40]=True
  close[floor_6,light_105]=True
  close[floor_6,floor_73]=True
  close[floor_6,floor_7]=True
  close[floor_6,wall_11]=True
  close[floor_6,wall_12]=True
  close[floor_6,wall_14]=True
  close[floor_6,wall_80]=True
  close[floor_6,mat_21]=True
  close[floor_6,light_62]=True
  close[floor_6,towel_rack_31]=True
  on[toy_314,filing_cabinet_305]=True
  close[controller_2054,table_281]=True
  close[towel_rack_31,floor_2]=True
  close[towel_rack_31,floor_3]=True
  close[towel_rack_31,floor_6]=True
  close[towel_rack_31,floor_73]=True
  close[towel_rack_31,floor_74]=True
  close[towel_rack_31,drawing_108]=True
  close[towel_rack_31,wall_12]=True
  close[towel_rack_31,wall_14]=True
  close[towel_rack_31,ceiling_15]=True
  close[towel_rack_31,wall_80]=True
  close[towel_rack_31,wall_81]=True
  close[towel_rack_31,ceiling_16]=True
  close[towel_rack_31,walllamp_25]=True
  close[towel_rack_31,ceiling_92]=True
  close[towel_rack_31,ceiling_93]=True
  close[towel_rack_31,light_62]=True
  facing[wall_76,drawing_108]=True
  on[fork_2004,desk_282]=True
  facing[bench_191,television_202]=True
  facing[bench_191,drawing_198]=True
  on[rag_2033,towel_rack_32]=True
  inside[tvstand_188,dining_room_163]=True
  close[wall_256,wall_260]=True
  close[wall_256,wall_261]=True
  close[wall_256,ceiling_267]=True
  close[wall_256,standingmirror_306]=True
  close[wall_256,window_275]=True
  close[wall_256,mat_308]=True
  close[wall_256,curtain_311]=True
  close[wall_256,curtain_312]=True
  close[wall_256,curtain_313]=True
  close[wall_256,floor_250]=True
  close[wall_256,couch_279]=True
  inside[drawing_198,dining_room_163]=True
  inside[curtain_111,bedroom_64]=True
  inside[curtain_111,curtain_112]=True
  close[bed_99,floor_65]=True
  close[bed_99,nightstand_98]=True
  close[bed_99,floor_67]=True
  close[bed_99,floor_66]=True
  close[bed_99,floor_68]=True
  close[bed_99,floor_70]=True
  close[bed_99,table_103]=True
  close[bed_99,sheets_2058]=True
  close[bed_99,mat_107]=True
  close[bed_99,wall_77]=True
  close[bed_99,wall_78]=True
  close[bed_99,curtain_111]=True
  close[bed_99,curtain_112]=True
  close[bed_99,pillow_113]=True
  close[bed_99,pillow_114]=True
  close[bed_99,vase_115]=True
  close[bed_99,window_84]=True
  close[bed_99,wall_79]=True
  close[bed_99,tablelamp_95]=True
  close[faucet_194,kitchen_counter_192]=True
  close[faucet_194,sink_193]=True
  close[faucet_194,cutting_board_228]=True
  close[faucet_194,floor_165]=True
  close[faucet_194,floor_164]=True
  close[faucet_194,toaster_231]=True
  close[faucet_194,floor_166]=True
  close[faucet_194,coffe_maker_236]=True
  close[faucet_194,wall_173]=True
  close[faucet_194,microwave_238]=True
  close[faucet_194,wall_174]=True
  close[faucet_194,ceiling_177]=True
  facing[floor_251,computer_321]=True
  facing[floor_251,drawing_307]=True
  facing[floor_251,drawing_309]=True
  facing[ceiling_181,drawing_197]=True
  facing[ceiling_181,drawing_198]=True
  inside[ground_coffee_2046,filing_cabinet_305]=True
  inside[ground_coffee_2046,home_office_246]=True
  inside[closetdrawer_146,bedroom_64]=True
  inside[closetdrawer_146,dresser_100]=True
  close[floor_7,chair_96]=True
  close[floor_7,shower_35]=True
  close[floor_7,wall_259]=True
  close[floor_7,toilet_37]=True
  close[floor_7,floor_6]=True
  close[floor_7,door_39]=True
  close[floor_7,floor_72]=True
  close[floor_7,floor_8]=True
  close[floor_7,light_105]=True
  close[floor_7,wall_11]=True
  close[floor_7,wall_10]=True
  close[floor_7,wall_82]=True
  close[floor_7,floor_247]=True
  close[floor_7,bookshelf_280]=True
  close[floor_7,walllamp_26]=True
  close[food_food_2055,table_189]=True
  facing[wall_259,drawing_307]=True
  facing[wall_259,drawing_309]=True
  close[food_jam_2013,cupboard_1000]=True
  close[stereo_2018,table_103]=True
  on[ceiling_182,wall_174]=True
  facing[chair_283,computer_321]=True
  close[ceiling_89,vase_115]=True
  close[ceiling_89,ceiling_86]=True
  close[ceiling_89,ceiling_88]=True
  close[ceiling_89,ceiling_90]=True
  close[ceiling_89,ceiling_92]=True
  close[ceiling_89,ceilinglamp_94]=True
  on[television_315,table_281]=True
  inside[pillow_114,bedroom_64]=True
  close[drawing_110,bookshelf_97]=True
  close[drawing_110,floor_69]=True
  close[drawing_110,drawing_198]=True
  close[drawing_110,doorjamb_104]=True
  close[drawing_110,floor_74]=True
  close[drawing_110,floor_170]=True
  close[drawing_110,wall_76]=True
  close[drawing_110,wall_175]=True
  close[drawing_110,wall_81]=True
  close[drawing_110,ceiling_180]=True
  close[drawing_110,door_183]=True
  close[drawing_110,ceiling_88]=True
  close[drawing_110,ceiling_93]=True
  close[ceiling_269,hanger_128]=True
  close[ceiling_269,hanger_129]=True
  close[ceiling_269,wall_258]=True
  close[ceiling_269,hanger_130]=True
  close[ceiling_269,wall_257]=True
  close[ceiling_269,wall_259]=True
  close[ceiling_269,hanger_131]=True
  close[ceiling_269,ceiling_264]=True
  close[ceiling_269,ceiling_268]=True
  close[ceiling_269,ceiling_270]=True
  close[ceiling_269,hanger_124]=True
  close[ceiling_269,doorjamb_273]=True
  close[ceiling_269,wall_83]=True
  close[ceiling_269,ceilinglamp_276]=True
  close[ceiling_269,bookshelf_280]=True
  close[ceiling_269,ceiling_91]=True
  close[ceiling_269,light_316]=True
  close[ceiling_269,hanger_125]=True
  close[ceiling_269,hanger_126]=True
  close[ceiling_269,hanger_127]=True
  inside[cup_1005,dining_room_163]=True
  close[drawing_309,wall_259]=True
  close[drawing_309,wall_262]=True
  close[drawing_309,ceiling_264]=True
  close[drawing_309,ceiling_265]=True
  close[drawing_309,filing_cabinet_305]=True
  close[drawing_309,walllamp_277]=True
  close[drawing_309,bookshelf_280]=True
  close[drawing_309,toy_314]=True
  on[couch_279,mat_308]=True
  on[couch_279,floor_255]=True
  inside[wall_78,bedroom_64]=True
  close[television_315,ceiling_268]=True
  close[television_315,ceilinglamp_276]=True
  close[television_315,mat_308]=True
  close[television_315,couch_279]=True
  close[television_315,floor_248]=True
  close[television_315,table_281]=True
  close[television_315,floor_250]=True
  close[television_315,floor_251]=True
  close[television_315,floor_254]=True
  on[oil_2053,table_189]=True
  close[cpuscreen_320,hanger_128]=True
  close[cpuscreen_320,wall_257]=True
  close[cpuscreen_320,hanger_130]=True
  close[cpuscreen_320,hanger_131]=True
  close[cpuscreen_320,hanger_132]=True
  close[cpuscreen_320,hanger_133]=True
  close[cpuscreen_320,hanger_129]=True
  close[cpuscreen_320,hanger_134]=True
  close[cpuscreen_320,wall_258]=True
  close[cpuscreen_320,closetdrawer_141]=True
  close[cpuscreen_320,closetdrawer_142]=True
  close[cpuscreen_320,closetdrawer_143]=True
  close[cpuscreen_320,closetdrawer_144]=True
  close[cpuscreen_320,ceiling_270]=True
  close[cpuscreen_320,closetdrawer_146]=True
  close[cpuscreen_320,closetdrawer_145]=True
  close[cpuscreen_320,desk_282]=True
  close[cpuscreen_320,chair_283]=True
  close[cpuscreen_320,light_316]=True
  close[cpuscreen_320,mouse_318]=True
  close[cpuscreen_320,mousepad_319]=True
  close[cpuscreen_320,computer_321]=True
  close[cpuscreen_320,keyboard_322]=True
  close[cpuscreen_320,floor_71]=True
  close[cpuscreen_320,wall_75]=True
  close[cpuscreen_320,wall_83]=True
  close[cpuscreen_320,ceiling_90]=True
  close[cpuscreen_320,dresser_100]=True
  close[cpuscreen_320,floor_253]=True
  close[cpuscreen_320,hanger_124]=True
  close[cpuscreen_320,hanger_125]=True
  close[cpuscreen_320,hanger_126]=True
  close[cpuscreen_320,hanger_127]=True
  close[floor_253,wall_257]=True
  close[floor_253,closetdrawer_141]=True
  close[floor_253,closetdrawer_142]=True
  close[floor_253,closetdrawer_143]=True
  close[floor_253,closetdrawer_144]=True
  close[floor_253,closetdrawer_145]=True
  close[floor_253,closetdrawer_146]=True
  close[floor_253,walllamp_278]=True
  close[floor_253,desk_282]=True
  close[floor_253,chair_283]=True
  close[floor_253,light_316]=True
  close[floor_253,powersocket_317]=True
  close[floor_253,mouse_318]=True
  close[floor_253,mousepad_319]=True
  close[floor_253,cpuscreen_320]=True
  close[floor_253,computer_321]=True
  close[floor_253,keyboard_322]=True
  close[floor_253,floor_71]=True
  close[floor_253,wall_75]=True
  close[floor_253,dresser_100]=True
  close[floor_253,floor_252]=True
  close[floor_253,floor_254]=True
  inside[food_jam_2013,cupboard_1000]=True
  inside[food_jam_2013,dining_room_163]=True
  close[floor_2,floor_3]=True
  close[floor_2,floor_4]=True
  close[floor_2,floor_6]=True
  close[floor_2,wall_9]=True
  close[floor_2,wall_12]=True
  close[floor_2,mat_21]=True
  close[floor_2,walllamp_25]=True
  close[floor_2,bathroom_counter_27]=True
  close[floor_2,sink_28]=True
  close[floor_2,faucet_29]=True
  close[floor_2,towel_rack_31]=True
  close[floor_2,floor_167]=True
  close[floor_2,door_39]=True
  close[floor_2,wall_176]=True
  close[floor_2,door_183]=True
  close[floor_2,light_62]=True
  close[floor_2,floor_74]=True
  close[floor_2,phone_205]=True
  close[floor_2,wall_81]=True
  close[floor_2,oven_229]=True
  close[floor_2,tray_230]=True
  facing[doorjamb_40,drawing_110]=True
  close[pencil_2050,table_103]=True
  inside[drawing_307,home_office_246]=True
  inside[ceiling_87,bedroom_64]=True
  on[sheets_2021,couch_279]=True
  close[chair_96,wall_258]=True
  close[chair_96,shower_35]=True
  close[chair_96,wall_259]=True
  close[chair_96,toilet_37]=True
  close[chair_96,floor_7]=True
  close[chair_96,floor_72]=True
  close[chair_96,wall_11]=True
  close[chair_96,doorjamb_273]=True
  close[chair_96,wall_82]=True
  close[chair_96,wall_83]=True
  close[chair_96,floor_252]=True
  close[chair_96,floor_247]=True
  close[chair_96,bookshelf_280]=True
  close[chair_96,ceiling_91]=True
  close[chair_96,light_316]=True
  close[chair_96,powersocket_317]=True
  facing[light_316,drawing_309]=True
  on[food_food_2009,table_103]=True
  close[bookshelf_195,drawing_197]=True
  close[bookshelf_195,drawing_198]=True
  close[bookshelf_195,floor_169]=True
  close[bookshelf_195,floor_170]=True
  close[bookshelf_195,wall_172]=True
  close[bookshelf_195,wall_175]=True
  close[bookshelf_195,ceiling_180]=True
  close[bookshelf_195,photoframe_219]=True
  close[bookshelf_195,check_2045]=True
  close[bookshelf_195,cutting_board_223]=True
  inside[ceiling_271,home_office_246]=True
  inside[purse_2022,home_office_246]=True
  inside[wall_81,bedroom_64]=True
  facing[floor_169,television_202]=True
  facing[floor_169,drawing_197]=True
  facing[floor_169,drawing_198]=True
  inside[novel_2042,home_office_246]=True
  inside[pillow_2006,dining_room_163]=True
  inside[ceiling_19,bathroom_1]=True
  inside[light_316,home_office_246]=True
  on[pillow_113,bed_99]=True
  on[television_202,tvstand_188]=True
  facing[ceiling_87,drawing_110]=True
  close[closetdrawer_143,hanger_128]=True
  close[closetdrawer_143,hanger_129]=True
  close[closetdrawer_143,hanger_130]=True
  close[closetdrawer_143,hanger_131]=True
  close[closetdrawer_143,hanger_132]=True
  close[closetdrawer_143,hanger_133]=True
  close[closetdrawer_143,hanger_134]=True
  close[closetdrawer_143,wall_257]=True
  close[closetdrawer_143,wall_258]=True
  close[closetdrawer_143,closetdrawer_141]=True
  close[closetdrawer_143,closetdrawer_142]=True
  close[closetdrawer_143,closetdrawer_144]=True
  close[closetdrawer_143,closetdrawer_145]=True
  close[closetdrawer_143,closetdrawer_146]=True
  close[closetdrawer_143,desk_282]=True
  close[closetdrawer_143,light_316]=True
  close[closetdrawer_143,powersocket_317]=True
  close[closetdrawer_143,mouse_318]=True
  close[closetdrawer_143,mousepad_319]=True
  close[closetdrawer_143,cpuscreen_320]=True
  close[closetdrawer_143,computer_321]=True
  close[closetdrawer_143,keyboard_322]=True
  close[closetdrawer_143,floor_71]=True
  close[closetdrawer_143,floor_72]=True
  close[closetdrawer_143,wall_75]=True
  close[closetdrawer_143,wall_83]=True
  close[closetdrawer_143,dresser_100]=True
  close[closetdrawer_143,floor_252]=True
  close[closetdrawer_143,floor_253]=True
  close[closetdrawer_143,hanger_124]=True
  close[closetdrawer_143,hanger_125]=True
  close[closetdrawer_143,hanger_126]=True
  close[closetdrawer_143,hanger_127]=True
  close[drawing_2014,filing_cabinet_305]=True
  facing[bed_99,drawing_109]=True
  facing[bed_99,drawing_110]=True
  close[food_food_2019,oven_229]=True
  inside[ceiling_264,home_office_246]=True
  close[cupboard_1000,blender_2048]=True
  close[cupboard_1000,bowl_1001]=True
  close[cupboard_1000,food_oatmeal_1002]=True
  close[cupboard_1000,fork_2035]=True
  close[cupboard_1000,food_jam_2013]=True
  inside[ceiling_90,bedroom_64]=True
  close[floor_166,floor_4]=True
  close[floor_166,wall_9]=True
  close[floor_166,mat_21]=True
  close[floor_166,walllamp_24]=True
  close[floor_166,bathroom_counter_27]=True
  close[floor_166,sink_28]=True
  close[floor_166,faucet_29]=True
  close[floor_166,floor_164]=True
  close[floor_166,floor_165]=True
  close[floor_166,floor_167]=True
  close[floor_166,wall_173]=True
  close[floor_166,wall_174]=True
  close[floor_166,table_189]=True
  close[floor_166,bench_191]=True
  close[floor_166,kitchen_counter_192]=True
  close[floor_166,sink_193]=True
  close[floor_166,faucet_194]=True
  close[floor_166,cutting_board_228]=True
  close[floor_166,oven_229]=True
  close[floor_166,tray_230]=True
  close[floor_166,freezer_234]=True
  close[floor_166,coffe_maker_236]=True
  close[floor_166,microwave_238]=True
  inside[hanger_126,bedroom_64]=True
  inside[hanger_126,dresser_100]=True
  close[wall_171,floor_168]=True
  close[wall_171,powersocket_201]=True
  close[wall_171,light_200]=True
  close[wall_171,television_202]=True
  close[wall_171,wall_172]=True
  close[wall_171,wall_173]=True
  close[wall_171,ceiling_178]=True
  close[wall_171,doorjamb_184]=True
  close[wall_171,maindoor_185]=True
  close[wall_171,tvstand_188]=True
  inside[clothes_shirt_2025,bedroom_64]=True
  inside[clothes_shirt_2025,dresser_100]=True
  inside[doorjamb_274,home_office_246]=True
  close[bench_191,mat_196]=True
  close[bench_191,floor_165]=True
  close[bench_191,floor_166]=True
  close[bench_191,floor_167]=True
  close[bench_191,floor_168]=True
  close[bench_191,orchid_199]=True
  close[bench_191,floor_164]=True
  close[bench_191,wall_173]=True
  close[bench_191,wall_174]=True
  close[bench_191,pillow_2006]=True
  close[bench_191,table_189]=True
  close[bench_191,bench_190]=True
  close[drawing_109,floor_65]=True
  close[drawing_109,floor_66]=True
  close[drawing_109,chair_101]=True
  close[drawing_109,wall_78]=True
  close[drawing_109,ceiling_85]=True
  close[mat_196,floor_167]=True
  close[mat_196,orchid_199]=True
  close[mat_196,floor_168]=True
  close[mat_196,wall_172]=True
  close[mat_196,wall_173]=True
  close[mat_196,wall_174]=True
  close[mat_196,wall_175]=True
  close[mat_196,table_189]=True
  close[mat_196,bench_190]=True
  close[mat_196,bench_191]=True
  facing[wall_77,drawing_109]=True
  on[faucet_29,bathroom_counter_27]=True
  inside[floor_74,bedroom_64]=True
  facing[television_202,drawing_197]=True
  inside[food_food_2009,bedroom_64]=True
  inside[shelf_38,bathroom_1]=True
  facing[floor_254,computer_321]=True
  inside[chair_283,home_office_246]=True
  inside[drawing_109,bedroom_64]=True
  inside[mousepad_319,home_office_246]=True
  facing[bookshelf_280,drawing_307]=True
  facing[bookshelf_280,drawing_309]=True
  on[check_2045,bookshelf_195]=True
  inside[wall_83,bedroom_64]=True
  close[ceiling_182,cutting_board_228]=True
  close[ceiling_182,bathroom_cabinet_36]=True
  close[ceiling_182,wall_9]=True
  close[ceiling_182,freezer_234]=True
  close[ceiling_182,stovefan_235]=True
  close[ceiling_182,coffe_maker_236]=True
  close[ceiling_182,wall_clock_204]=True
  close[ceiling_182,wall_174]=True
  close[ceiling_182,microwave_238]=True
  close[ceiling_182,wall_173]=True
  close[ceiling_182,ceiling_177]=True
  close[ceiling_182,ceiling_20]=True
  close[ceiling_182,ceiling_181]=True
  close[ceiling_182,walllamp_24]=True
  close[ceiling_182,ceilinglamp_187]=True
  close[ceiling_182,faucet_29]=True
  close[ceilinglamp_186,wall_172]=True
  close[ceilinglamp_186,wall_175]=True
  close[ceilinglamp_186,ceiling_178]=True
  close[ceilinglamp_186,ceiling_179]=True
  close[ceilinglamp_186,ceiling_180]=True
  close[ceilinglamp_186,ceiling_181]=True
  inside[stereo_2018,bedroom_64]=True
  inside[ceiling_267,home_office_246]=True
  on[ceiling_18,wall_10]=True
  inside[ceiling_93,bedroom_64]=True
  between[door_183,bedroom_64]=True
  between[door_183,dining_room_163]=True
  on[bookshelf_280,floor_247]=True
  facing[wall_258,drawing_309]=True
  close[tray_230,kitchen_counter_192]=True
  close[tray_230,floor_2]=True
  close[tray_230,floor_3]=True
  close[tray_230,bathroom_cabinet_36]=True
  close[tray_230,oven_229]=True
  close[tray_230,floor_166]=True
  close[tray_230,floor_4]=True
  close[tray_230,floor_167]=True
  close[tray_230,wall_9]=True
  close[tray_230,freezer_234]=True
  close[tray_230,stovefan_235]=True
  close[tray_230,wall_12]=True
  close[tray_230,wall_174]=True
  close[tray_230,wall_176]=True
  close[tray_230,mat_21]=True
  close[tray_230,walllamp_24]=True
  close[tray_230,bathroom_counter_27]=True
  close[tray_230,sink_28]=True
  close[tray_230,faucet_29]=True
  inside[video_game_controller_2028,bedroom_64]=True
  close[freezer_234,food_food_2052]=True
  close[freezer_234,wall_9]=True
  close[freezer_234,walllamp_24]=True
  close[freezer_234,floor_164]=True
  close[freezer_234,floor_165]=True
  close[freezer_234,floor_166]=True
  close[freezer_234,wall_173]=True
  close[freezer_234,wall_174]=True
  close[freezer_234,ceiling_182]=True
  close[freezer_234,table_189]=True
  close[freezer_234,kitchen_counter_192]=True
  close[freezer_234,food_food_2015]=True
  close[freezer_234,cutting_board_228]=True
  close[freezer_234,oven_229]=True
  close[freezer_234,tray_230]=True
  close[freezer_234,stovefan_235]=True
  close[freezer_234,coffe_maker_236]=True
  close[freezer_234,milk_1003]=True
  close[freezer_234,microwave_238]=True
  close[freezer_234,ground_coffee_1004]=True
  close[freezer_234,cup_1005]=True
  close[freezer_234,juice_1006]=True
  close[freezer_234,juice_2043]=True
  close[floor_255,wall_261]=True
  close[floor_255,mat_308]=True
  close[floor_255,pillow_310]=True
  close[floor_255,couch_279]=True
  close[floor_255,table_281]=True
  close[floor_255,floor_250]=True
  close[floor_255,floor_254]=True
  inside[floor_251,home_office_246]=True
  facing[pillow_310,television_315]=True
  inside[curtain_312,home_office_246]=True
  inside[curtain_312,curtain_311]=True
  facing[floor_164,wall_clock_204]=True
  close[piano_bench_2005,floor_254]=True
  inside[floor_5,bathroom_1]=True
  inside[oil_2053,dining_room_163]=True
  close[clothes_skirt_2010,couch_279]=True
  close[food_carrot_2016,kitchen_counter_192]=True
  facing[tvstand_188,television_202]=True
  facing[tvstand_188,drawing_197]=True
  facing[tvstand_188,drawing_198]=True
  inside[ceilinglamp_276,home_office_246]=True
  on[novel_2034,table_189]=True
  inside[hanger_102,bedroom_64]=True
  on[food_rice_2038,kitchen_counter_192]=True
  close[wall_261,wall_256]=True
  close[wall_261,wall_263]=True
  close[wall_261,ceiling_267]=True
  close[wall_261,ceiling_271]=True
  close[wall_261,ceiling_272]=True
  close[wall_261,doorjamb_274]=True
  close[wall_261,window_275]=True
  close[wall_261,mat_308]=True
  close[wall_261,pillow_310]=True
  close[wall_261,couch_279]=True
  close[wall_261,curtain_312]=True
  close[wall_261,table_281]=True
  close[wall_261,floor_250]=True
  close[wall_261,curtain_311]=True
  close[wall_261,floor_254]=True
  close[wall_261,floor_255]=True
  inside[centerpiece_2037,filing_cabinet_305]=True
  inside[centerpiece_2037,home_office_246]=True
  facing[floor_65,drawing_109]=True
  close[drawing_307,hanger_289]=True
  close[drawing_307,hanger_291]=True
  close[drawing_307,wall_260]=True
  close[drawing_307,hanger_293]=True
  close[drawing_307,wall_262]=True
  close[drawing_307,closetdrawer_296]=True
  close[drawing_307,ceiling_265]=True
  close[drawing_307,ceiling_266]=True
  close[drawing_307,closetdrawer_301]=True
  close[drawing_307,filing_cabinet_305]=True
  close[drawing_307,walllamp_277]=True
  close[drawing_307,toy_314]=True
  close[drawing_307,dresser_284]=True
  close[drawing_307,hanger_285]=True
  close[curtain_312,wall_256]=True
  close[curtain_312,wall_261]=True
  close[curtain_312,ceiling_267]=True
  close[curtain_312,ceiling_272]=True
  close[curtain_312,window_275]=True
  close[curtain_312,mat_308]=True
  close[curtain_312,couch_279]=True
  close[curtain_312,curtain_313]=True
  close[curtain_312,floor_250]=True
  close[curtain_312,curtain_311]=True
  inside[wall_14,bathroom_1]=True
  on[closetdrawer_144,closetdrawer_146]=True
  inside[sheets_2062,filing_cabinet_305]=True
  inside[sheets_2062,home_office_246]=True
  inside[wallshelf_34,bathroom_1]=True
  facing[powersocket_317,drawing_309]=True
  close[ceiling_17,shower_35]=True
  close[ceiling_17,wall_259]=True
  close[ceiling_17,ceiling_264]=True
  close[ceiling_17,light_105]=True
  close[ceiling_17,wall_10]=True
  close[ceiling_17,wall_11]=True
  close[ceiling_17,ceiling_16]=True
  close[ceiling_17,wall_82]=True
  close[ceiling_17,ceiling_18]=True
  close[ceiling_17,ceilinglamp_23]=True
  close[ceiling_17,walllamp_26]=True
  close[ceiling_17,ceiling_91]=True
  close[toilet_37,chair_96]=True
  close[toilet_37,wall_258]=True
  close[toilet_37,shower_35]=True
  close[toilet_37,wall_259]=True
  close[toilet_37,floor_7]=True
  close[toilet_37,floor_72]=True
  close[toilet_37,wall_11]=True
  close[toilet_37,wall_82]=True
  close[toilet_37,wall_83]=True
  close[toilet_37,floor_247]=True
  close[toilet_37,bookshelf_280]=True
  close[toilet_37,floor_252]=True
  inside[floor_254,home_office_246]=True
  inside[hanger_295,dresser_284]=True
  inside[hanger_295,home_office_246]=True
  close[form_2029,bookshelf_97]=True
  facing[cutting_board_223,drawing_108]=True
  close[ceiling_88,bookshelf_97]=True
  close[ceiling_88,drawing_198]=True
  close[ceiling_88,wall_76]=True
  close[ceiling_88,drawing_110]=True
  close[ceiling_88,wall_79]=True
  close[ceiling_88,wall_81]=True
  close[ceiling_88,ceiling_87]=True
  close[ceiling_88,ceiling_89]=True
  close[ceiling_88,ceiling_93]=True
  close[ceiling_88,ceilinglamp_94]=True
  inside[television_202,dining_room_163]=True
  close[wall_263,wall_257]=True
  close[wall_263,wall_261]=True
  close[wall_263,ceiling_271]=True
  close[wall_263,doorjamb_274]=True
  close[wall_263,mat_308]=True
  close[wall_263,walllamp_278]=True
  close[wall_263,couch_279]=True
  close[wall_263,chair_283]=True
  close[wall_263,floor_254]=True
  inside[floor_69,bedroom_64]=True
  close[ceiling_268,ceiling_265]=True
  close[ceiling_268,ceiling_267]=True
  close[ceiling_268,ceiling_269]=True
  close[ceiling_268,ceiling_271]=True
  close[ceiling_268,ceilinglamp_276]=True
  close[ceiling_268,television_315]=True
  inside[juice_1006,freezer_234]=True
  inside[juice_1006,dining_room_163]=True
  facing[floor_247,drawing_307]=True
  facing[floor_247,drawing_309]=True
  facing[floor_74,drawing_108]=True
  facing[floor_74,drawing_110]=True
  on[bench_191,floor_167]=True
  inside[floor_166,dining_room_163]=True
  inside[cupboard_1000,dining_room_163]=True
  inside[ceiling_17,bathroom_1]=True
  on[ceiling_179,wall_172]=True
  facing[nightstand_98,drawing_110]=True
  close[floor_252,wall_257]=True
  close[floor_252,wall_258]=True
  close[floor_252,wall_259]=True
  close[floor_252,closetdrawer_143]=True
  close[floor_252,closetdrawer_144]=True
  close[floor_252,doorjamb_273]=True
  close[floor_252,closetdrawer_146]=True
  close[floor_252,bookshelf_280]=True
  close[floor_252,desk_282]=True
  close[floor_252,toilet_37]=True
  close[floor_252,light_316]=True
  close[floor_252,powersocket_317]=True
  close[floor_252,mouse_318]=True
  close[floor_252,mousepad_319]=True
  close[floor_252,computer_321]=True
  close[floor_252,floor_72]=True
  close[floor_252,wall_83]=True
  close[floor_252,chair_96]=True
  close[floor_252,floor_247]=True
  close[floor_252,floor_251]=True
  close[floor_252,floor_253]=True
  on[closetdrawer_143,closetdrawer_144]=True
  inside[broom_2049,dining_room_163]=True
  facing[wall_176,drawing_198]=True
  inside[wall_262,home_office_246]=True
  inside[wall_175,dining_room_163]=True
  close[wall_258,hanger_128]=True
  close[wall_258,hanger_129]=True
  close[wall_258,hanger_130]=True
  close[wall_258,hanger_131]=True
  close[wall_258,wall_257]=True
  close[wall_258,wall_259]=True
  close[wall_258,wall_11]=True
  close[wall_258,ceiling_269]=True
  close[wall_258,closetdrawer_143]=True
  close[wall_258,closetdrawer_144]=True
  close[wall_258,doorjamb_273]=True
  close[wall_258,closetdrawer_146]=True
  close[wall_258,bookshelf_280]=True
  close[wall_258,desk_282]=True
  close[wall_258,shower_35]=True
  close[wall_258,toilet_37]=True
  close[wall_258,light_316]=True
  close[wall_258,powersocket_317]=True
  close[wall_258,mouse_318]=True
  close[wall_258,mousepad_319]=True
  close[wall_258,cpuscreen_320]=True
  close[wall_258,computer_321]=True
  close[wall_258,keyboard_322]=True
  close[wall_258,floor_72]=True
  close[wall_258,wall_75]=True
  close[wall_258,wall_82]=True
  close[wall_258,wall_83]=True
  close[wall_258,ceiling_91]=True
  close[wall_258,chair_96]=True
  close[wall_258,dresser_100]=True
  close[wall_258,hanger_124]=True
  close[wall_258,floor_252]=True
  close[wall_258,hanger_125]=True
  close[wall_258,hanger_126]=True
  close[wall_258,hanger_127]=True
  close[chair_101,floor_65]=True
  close[chair_101,floor_66]=True
  close[chair_101,floor_67]=True
  close[chair_101,mat_107]=True
  close[chair_101,drawing_109]=True
  close[chair_101,wall_78]=True
  close[chair_101,wall_77]=True
  close[chair_101,ceiling_85]=True
  on[clothes_skirt_2010,couch_279]=True
  close[mat_107,floor_65]=True
  close[mat_107,floor_66]=True
  close[mat_107,floor_67]=True
  close[mat_107,floor_68]=True
  close[mat_107,floor_69]=True
  close[mat_107,floor_70]=True
  close[mat_107,floor_71]=True
  close[mat_107,wall_77]=True
  close[mat_107,wall_78]=True
  close[mat_107,wall_79]=True
  close[mat_107,window_84]=True
  close[mat_107,tablelamp_95]=True
  close[mat_107,nightstand_98]=True
  close[mat_107,bed_99]=True
  close[mat_107,chair_101]=True
  close[mat_107,table_103]=True
  close[mat_107,curtain_111]=True
  close[mat_107,curtain_112]=True
  close[mat_107,pillow_113]=True
  close[mat_107,pillow_114]=True
  close[mat_107,vase_115]=True
  inside[floor_169,dining_room_163]=True
  facing[ceiling_182,wall_clock_204]=True
  close[standingmirror_306,wall_256]=True
  close[standingmirror_306,wall_260]=True
  close[standingmirror_306,floor_249]=True
  close[standingmirror_306,hanger_295]=True
  close[standingmirror_306,closetdrawer_296]=True
  close[standingmirror_306,ceiling_266]=True
  close[standingmirror_306,closetdrawer_299]=True
  close[standingmirror_306,ceiling_267]=True
  close[standingmirror_306,window_275]=True
  close[standingmirror_306,curtain_313]=True
  close[standingmirror_306,floor_250]=True
  close[standingmirror_306,dresser_284]=True
  close[standingmirror_306,hanger_287]=True
  inside[wall_10,bathroom_1]=True
  facing[table_281,computer_321]=True
  facing[table_281,television_315]=True
  facing[table_281,drawing_307]=True
  facing[table_281,drawing_309]=True
  inside[sheets_2058,bedroom_64]=True
  inside[hanger_133,bedroom_64]=True
  inside[hanger_133,dresser_100]=True
  on[pillow_114,bed_99]=True
  inside[tray_230,dining_room_163]=True
  inside[tray_230,oven_229]=True
  facing[wall_175,drawing_108]=True
  facing[wall_175,drawing_197]=True
  facing[wall_175,drawing_198]=True
  on[food_food_2055,table_189]=True
  inside[ceiling_178,dining_room_163]=True
  close[table_103,stereo_2018]=True
  close[table_103,bed_99]=True
  close[table_103,floor_67]=True
  close[table_103,floor_69]=True
  close[table_103,floor_70]=True
  close[table_103,floor_71]=True
  close[table_103,pencil_2050]=True
  close[table_103,floor_73]=True
  close[table_103,mat_107]=True
  close[table_103,video_game_controller_2028]=True
  close[table_103,vase_115]=True
  close[table_103,food_food_2009]=True
  facing[stovefan_235,wall_clock_204]=True
  close[drawing_108,door_39]=True
  close[drawing_108,doorjamb_40]=True
  close[drawing_108,floor_74]=True
  close[drawing_108,wall_12]=True
  close[drawing_108,phone_205]=True
  close[drawing_108,wall_14]=True
  close[drawing_108,ceiling_15]=True
  close[drawing_108,wall_80]=True
  close[drawing_108,wall_81]=True
  close[drawing_108,ceiling_16]=True
  close[drawing_108,walllamp_25]=True
  close[drawing_108,ceiling_92]=True
  close[drawing_108,ceiling_93]=True
  close[drawing_108,light_62]=True
  close[drawing_108,towel_rack_31]=True
  inside[closetdrawer_142,bedroom_64]=True
  inside[closetdrawer_142,dresser_100]=True
  facing[wall_78,drawing_109]=True
  close[powersocket_201,floor_164]=True
  close[powersocket_201,floor_165]=True
  close[powersocket_201,light_200]=True
  close[powersocket_201,floor_168]=True
  close[powersocket_201,wall_171]=True
  close[powersocket_201,wall_173]=True
  close[powersocket_201,doorjamb_184]=True
  close[powersocket_201,maindoor_185]=True
  facing[floor_165,wall_clock_204]=True
  inside_char[char,bedroom_64]=True
  facing[table_189,drawing_197]=True
  facing[table_189,drawing_198]=True
  facing[toy_314,drawing_307]=True
  on[towel_2011,kitchen_counter_192]=True
  close[hanger_129,hanger_128]=True
  close[hanger_129,wall_257]=True
  close[hanger_129,hanger_130]=True
  close[hanger_129,hanger_131]=True
  close[hanger_129,hanger_132]=True
  close[hanger_129,hanger_133]=True
  close[hanger_129,hanger_134]=True
  close[hanger_129,wall_258]=True
  close[hanger_129,closetdrawer_141]=True
  close[hanger_129,ceiling_270]=True
  close[hanger_129,closetdrawer_143]=True
  close[hanger_129,closetdrawer_144]=True
  close[hanger_129,doorjamb_273]=True
  close[hanger_129,ceiling_269]=True
  close[hanger_129,desk_282]=True
  close[hanger_129,light_316]=True
  close[hanger_129,mouse_318]=True
  close[hanger_129,mousepad_319]=True
  close[hanger_129,cpuscreen_320]=True
  close[hanger_129,keyboard_322]=True
  close[hanger_129,wall_75]=True
  close[hanger_129,wall_83]=True
  close[hanger_129,ceiling_90]=True
  close[hanger_129,ceiling_91]=True
  close[hanger_129,dresser_100]=True
  close[hanger_129,hanger_124]=True
  close[hanger_129,hanger_125]=True
  close[hanger_129,hanger_126]=True
  close[hanger_129,hanger_127]=True
  close[cup_2008,kitchen_counter_192]=True
  facing[ceiling_267,television_315]=True
  facing[ceiling_267,drawing_307]=True
  inside[drawing_197,dining_room_163]=True
  close[nightstand_98,floor_67]=True
  close[nightstand_98,floor_68]=True
  close[nightstand_98,bed_99]=True
  close[nightstand_98,mat_107]=True
  close[nightstand_98,wall_77]=True
  close[nightstand_98,curtain_111]=True
  close[nightstand_98,curtain_112]=True
  close[nightstand_98,pillow_113]=True
  close[nightstand_98,wall_79]=True
  close[nightstand_98,pillow_114]=True
  close[nightstand_98,window_84]=True
  close[nightstand_98,tablelamp_95]=True
  inside[doorjamb_104,bedroom_64]=True
  inside[closetdrawer_145,bedroom_64]=True
  inside[closetdrawer_145,dresser_100]=True
  inside[ceiling_181,dining_room_163]=True
  inside[hanger_129,bedroom_64]=True
  inside[hanger_129,dresser_100]=True
  close[wall_9,floor_2]=True
  close[wall_9,floor_3]=True
  close[wall_9,floor_4]=True
  close[wall_9,floor_5]=True
  close[wall_9,wall_12]=True
  close[wall_9,wall_13]=True
  close[wall_9,ceiling_15]=True
  close[wall_9,ceiling_19]=True
  close[wall_9,ceiling_20]=True
  close[wall_9,mat_21]=True
  close[wall_9,curtain_22]=True
  close[wall_9,ceilinglamp_23]=True
  close[wall_9,walllamp_24]=True
  close[wall_9,bathroom_counter_27]=True
  close[wall_9,sink_28]=True
  close[wall_9,faucet_29]=True
  close[wall_9,towel_rack_33]=True
  close[wall_9,wallshelf_34]=True
  close[wall_9,bathroom_cabinet_36]=True
  close[wall_9,floor_166]=True
  close[wall_9,wall_174]=True
  close[wall_9,wall_176]=True
  close[wall_9,ceiling_182]=True
  close[wall_9,window_61]=True
  close[wall_9,wall_clock_204]=True
  close[wall_9,oven_229]=True
  close[wall_9,tray_230]=True
  close[wall_9,freezer_234]=True
  close[wall_9,stovefan_235]=True
  close[food_salt_2057,sink_28]=True
  close[fork_2004,desk_282]=True
  inside[pillow_113,bedroom_64]=True
  close[doorjamb_40,floor_6]=True
  close[doorjamb_40,door_39]=True
  close[doorjamb_40,light_105]=True
  close[doorjamb_40,floor_73]=True
  close[doorjamb_40,wall_11]=True
  close[doorjamb_40,drawing_108]=True
  close[doorjamb_40,wall_12]=True
  close[doorjamb_40,wall_14]=True
  close[doorjamb_40,wall_80]=True
  close[doorjamb_40,ceiling_16]=True
  close[doorjamb_40,wall_82]=True
  close[doorjamb_40,wall_81]=True
  close[doorjamb_40,ceiling_92]=True
  close[doorjamb_40,light_62]=True
  facing[ceilinglamp_276,computer_321]=True
  facing[ceilinglamp_276,drawing_307]=True
  facing[ceilinglamp_276,drawing_309]=True
  inside[bench_190,dining_room_163]=True
  close[wall_173,floor_164]=True
  close[wall_173,floor_165]=True
  close[wall_173,floor_166]=True
  close[wall_173,floor_168]=True
  close[wall_173,wall_171]=True
  close[wall_173,wall_174]=True
  close[wall_173,ceiling_177]=True
  close[wall_173,ceiling_178]=True
  close[wall_173,ceiling_182]=True
  close[wall_173,doorjamb_184]=True
  close[wall_173,maindoor_185]=True
  close[wall_173,ceilinglamp_187]=True
  close[wall_173,table_189]=True
  close[wall_173,bench_191]=True
  close[wall_173,kitchen_counter_192]=True
  close[wall_173,sink_193]=True
  close[wall_173,faucet_194]=True
  close[wall_173,mat_196]=True
  close[wall_173,orchid_199]=True
  close[wall_173,light_200]=True
  close[wall_173,powersocket_201]=True
  close[wall_173,cutting_board_228]=True
  close[wall_173,toaster_231]=True
  close[wall_173,freezer_234]=True
  close[wall_173,coffe_maker_236]=True
  close[wall_173,microwave_238]=True
  close[wall_260,wall_256]=True
  close[wall_260,wall_262]=True
  close[wall_260,ceiling_265]=True
  close[wall_260,ceiling_266]=True
  close[wall_260,ceiling_267]=True
  close[wall_260,window_275]=True
  close[wall_260,dresser_284]=True
  close[wall_260,hanger_285]=True
  close[wall_260,hanger_287]=True
  close[wall_260,hanger_289]=True
  close[wall_260,hanger_291]=True
  close[wall_260,hanger_293]=True
  close[wall_260,hanger_295]=True
  close[wall_260,closetdrawer_296]=True
  close[wall_260,closetdrawer_299]=True
  close[wall_260,closetdrawer_301]=True
  close[wall_260,standingmirror_306]=True
  close[wall_260,drawing_307]=True
  close[wall_260,curtain_313]=True
  close[wall_260,floor_248]=True
  close[wall_260,floor_249]=True
  close[wall_260,floor_250]=True
  close[window_275,wall_256]=True
  close[window_275,wall_260]=True
  close[window_275,wall_261]=True
  close[window_275,ceiling_267]=True
  close[window_275,standingmirror_306]=True
  close[window_275,mat_308]=True
  close[window_275,curtain_311]=True
  close[window_275,curtain_312]=True
  close[window_275,curtain_313]=True
  close[window_275,floor_250]=True
  close[window_275,couch_279]=True
  facing[curtain_312,television_315]=True
  inside[bookshelf_97,bedroom_64]=True
  close[photoframe_219,bookshelf_195]=True
  close[photoframe_219,drawing_197]=True
  close[photoframe_219,floor_169]=True
  close[photoframe_219,television_202]=True
  close[photoframe_219,wall_172]=True
  close[photoframe_219,tvstand_188]=True
  inside[wall_clock_2032,bathroom_1]=True
  facing[ceiling_177,wall_clock_204]=True
  inside[window_61,bathroom_1]=True
  on[piano_bench_2047,floor_254]=True
  close[wall_11,wall_258]=True
  close[wall_11,wall_259]=True
  close[wall_11,floor_6]=True
  close[wall_11,floor_7]=True
  close[wall_11,floor_8]=True
  close[wall_11,ceiling_264]=True
  close[wall_11,wall_10]=True
  close[wall_11,wall_14]=True
  close[wall_11,ceiling_16]=True
  close[wall_11,ceiling_17]=True
  close[wall_11,doorjamb_273]=True
  close[wall_11,ceiling_18]=True
  close[wall_11,ceilinglamp_23]=True
  close[wall_11,bookshelf_280]=True
  close[wall_11,walllamp_26]=True
  close[wall_11,shower_35]=True
  close[wall_11,toilet_37]=True
  close[wall_11,door_39]=True
  close[wall_11,doorjamb_40]=True
  close[wall_11,floor_72]=True
  close[wall_11,wall_80]=True
  close[wall_11,wall_82]=True
  close[wall_11,wall_83]=True
  close[wall_11,ceiling_91]=True
  close[wall_11,chair_96]=True
  close[wall_11,light_105]=True
  close[wall_11,floor_247]=True
  close[blow_dryer_2059,bathroom_counter_27]=True
  facing[floor_71,drawing_109]=True
  close[ceiling_16,doorjamb_40]=True
  close[ceiling_16,light_105]=True
  close[ceiling_16,wall_11]=True
  close[ceiling_16,drawing_108]=True
  close[ceiling_16,wall_12]=True
  close[ceiling_16,wall_14]=True
  close[ceiling_16,ceiling_15]=True
  close[ceiling_16,wall_80]=True
  close[ceiling_16,ceiling_17]=True
  close[ceiling_16,ceiling_19]=True
  close[ceiling_16,ceilinglamp_23]=True
  close[ceiling_16,ceiling_92]=True
  close[ceiling_16,light_62]=True
  close[ceiling_16,towel_rack_31]=True
  inside[standingmirror_306,home_office_246]=True
  close[bathroom_cabinet_36,oven_229]=True
  close[bathroom_cabinet_36,tray_230]=True
  close[bathroom_cabinet_36,wall_9]=True
  close[bathroom_cabinet_36,stovefan_235]=True
  close[bathroom_cabinet_36,wall_clock_204]=True
  close[bathroom_cabinet_36,wall_12]=True
  close[bathroom_cabinet_36,wall_174]=True
  close[bathroom_cabinet_36,ceiling_15]=True
  close[bathroom_cabinet_36,wall_176]=True
  close[bathroom_cabinet_36,phone_205]=True
  close[bathroom_cabinet_36,ceiling_20]=True
  close[bathroom_cabinet_36,ceiling_181]=True
  close[bathroom_cabinet_36,ceiling_182]=True
  close[bathroom_cabinet_36,walllamp_24]=True
  close[bathroom_cabinet_36,walllamp_25]=True
  close[bathroom_cabinet_36,bathroom_counter_27]=True
  close[bathroom_cabinet_36,sink_28]=True
  close[bathroom_cabinet_36,faucet_29]=True
  on[stamp_2056,bookshelf_280]=True
  surfaces[floor_2] = True
  surfaces[floor_3] = True
  surfaces[floor_4] = True
  surfaces[floor_5] = True
  surfaces[floor_6] = True
  surfaces[floor_7] = True
  surfaces[floor_8] = True
  sittable[mat_21] = True
  grabbable[mat_21] = True
  movable[mat_21] = True
  lieable[mat_21] = True
  surfaces[mat_21] = True
  movable[curtain_22] = True
  can_open[curtain_22] = True
  cover_object[curtain_22] = True
  surfaces[bathroom_counter_27] = True
  recipient[sink_28] = True
  containers[sink_28] = True
  has_switch[faucet_29] = True
  lieable[bathtub_30] = True
  sittable[bathtub_30] = True
  grabbable[towel_rack_31] = True
  movable[towel_rack_31] = True
  surfaces[towel_rack_31] = True
  grabbable[towel_rack_32] = True
  movable[towel_rack_32] = True
  surfaces[towel_rack_32] = True
  grabbable[towel_rack_33] = True
  movable[towel_rack_33] = True
  surfaces[towel_rack_33] = True
  can_open[bathroom_cabinet_36] = True
  surfaces[bathroom_cabinet_36] = True
  containers[bathroom_cabinet_36] = True
  can_open[toilet_37] = True
  containers[toilet_37] = True
  sittable[toilet_37] = True
  can_open[door_39] = True
  has_switch[light_62] = True
  has_plug[light_62] = True
  surfaces[floor_65] = True
  surfaces[floor_66] = True
  surfaces[floor_67] = True
  surfaces[floor_68] = True
  surfaces[floor_69] = True
  surfaces[floor_70] = True
  surfaces[floor_71] = True
  surfaces[floor_72] = True
  surfaces[floor_73] = True
  surfaces[floor_74] = True
  has_switch[tablelamp_95] = True
  grabbable[chair_96] = True
  movable[chair_96] = True
  surfaces[chair_96] = True
  sittable[chair_96] = True
  can_open[bookshelf_97] = True
  surfaces[bookshelf_97] = True
  containers[bookshelf_97] = True
  can_open[nightstand_98] = True
  surfaces[nightstand_98] = True
  containers[nightstand_98] = True
  lieable[bed_99] = True
  surfaces[bed_99] = True
  sittable[bed_99] = True
  can_open[dresser_100] = True
  containers[dresser_100] = True
  grabbable[chair_101] = True
  movable[chair_101] = True
  surfaces[chair_101] = True
  sittable[chair_101] = True
  grabbable[hanger_102] = True
  movable[hanger_102] = True
  hangable[hanger_102] = True
  movable[table_103] = True
  surfaces[table_103] = True
  has_switch[light_105] = True
  has_plug[light_105] = True
  sittable[mat_107] = True
  grabbable[mat_107] = True
  movable[mat_107] = True
  lieable[mat_107] = True
  surfaces[mat_107] = True
  has_paper[drawing_108] = True
  cuttable[drawing_108] = True
  grabbable[drawing_108] = True
  movable[drawing_108] = True
  lookable[drawing_108] = True
  has_paper[drawing_109] = True
  cuttable[drawing_109] = True
  grabbable[drawing_109] = True
  movable[drawing_109] = True
  lookable[drawing_109] = True
  has_paper[drawing_110] = True
  cuttable[drawing_110] = True
  grabbable[drawing_110] = True
  movable[drawing_110] = True
  lookable[drawing_110] = True
  movable[curtain_111] = True
  can_open[curtain_111] = True
  cover_object[curtain_111] = True
  movable[curtain_112] = True
  can_open[curtain_112] = True
  cover_object[curtain_112] = True
  grabbable[pillow_113] = True
  movable[pillow_113] = True
  grabbable[pillow_114] = True
  movable[pillow_114] = True
  grabbable[hanger_124] = True
  movable[hanger_124] = True
  hangable[hanger_124] = True
  grabbable[hanger_125] = True
  movable[hanger_125] = True
  hangable[hanger_125] = True
  grabbable[hanger_126] = True
  movable[hanger_126] = True
  hangable[hanger_126] = True
  grabbable[hanger_127] = True
  movable[hanger_127] = True
  hangable[hanger_127] = True
  grabbable[hanger_128] = True
  movable[hanger_128] = True
  hangable[hanger_128] = True
  grabbable[hanger_129] = True
  movable[hanger_129] = True
  hangable[hanger_129] = True
  grabbable[hanger_130] = True
  movable[hanger_130] = True
  hangable[hanger_130] = True
  grabbable[hanger_131] = True
  movable[hanger_131] = True
  hangable[hanger_131] = True
  grabbable[hanger_132] = True
  movable[hanger_132] = True
  hangable[hanger_132] = True
  grabbable[hanger_133] = True
  movable[hanger_133] = True
  hangable[hanger_133] = True
  grabbable[hanger_134] = True
  movable[hanger_134] = True
  hangable[hanger_134] = True
  surfaces[floor_164] = True
  surfaces[floor_165] = True
  surfaces[floor_166] = True
  surfaces[floor_167] = True
  surfaces[floor_168] = True
  surfaces[floor_169] = True
  surfaces[floor_170] = True
  can_open[door_183] = True
  surfaces[tvstand_188] = True
  movable[table_189] = True
  surfaces[table_189] = True
  movable[bench_190] = True
  lieable[bench_190] = True
  surfaces[bench_190] = True
  sittable[bench_190] = True
  movable[bench_191] = True
  lieable[bench_191] = True
  surfaces[bench_191] = True
  sittable[bench_191] = True
  surfaces[kitchen_counter_192] = True
  recipient[sink_193] = True
  containers[sink_193] = True
  has_switch[faucet_194] = True
  can_open[bookshelf_195] = True
  surfaces[bookshelf_195] = True
  containers[bookshelf_195] = True
  sittable[mat_196] = True
  grabbable[mat_196] = True
  movable[mat_196] = True
  lieable[mat_196] = True
  surfaces[mat_196] = True
  has_paper[drawing_197] = True
  cuttable[drawing_197] = True
  grabbable[drawing_197] = True
  movable[drawing_197] = True
  lookable[drawing_197] = True
  has_paper[drawing_198] = True
  cuttable[drawing_198] = True
  grabbable[drawing_198] = True
  movable[drawing_198] = True
  lookable[drawing_198] = True
  has_switch[light_200] = True
  has_plug[light_200] = True
  has_switch[television_202] = True
  lookable[television_202] = True
  has_plug[television_202] = True
  grabbable[wall_clock_204] = True
  movable[wall_clock_204] = True
  has_plug[wall_clock_204] = True
  lookable[wall_clock_204] = True
  has_switch[wall_clock_204] = True
  grabbable[phone_205] = True
  movable[phone_205] = True
  has_switch[phone_205] = True
  has_plug[phone_205] = True
  grabbable[cutting_board_223] = True
  movable[cutting_board_223] = True
  surfaces[cutting_board_223] = True
  grabbable[cutting_board_228] = True
  movable[cutting_board_228] = True
  surfaces[cutting_board_228] = True
  has_plug[oven_229] = True
  can_open[oven_229] = True
  containers[oven_229] = True
  has_switch[oven_229] = True
  grabbable[tray_230] = True
  movable[tray_230] = True
  surfaces[tray_230] = True
  movable[toaster_231] = True
  has_switch[toaster_231] = True
  has_plug[toaster_231] = True
  has_plug[freezer_234] = True
  can_open[freezer_234] = True
  containers[freezer_234] = True
  has_switch[freezer_234] = True
  containers[coffe_maker_236] = True
  movable[coffe_maker_236] = True
  recipient[coffe_maker_236] = True
  has_plug[coffe_maker_236] = True
  can_open[coffe_maker_236] = True
  has_switch[coffe_maker_236] = True
  has_plug[microwave_238] = True
  can_open[microwave_238] = True
  containers[microwave_238] = True
  has_switch[microwave_238] = True
  surfaces[floor_247] = True
  surfaces[floor_248] = True
  surfaces[floor_249] = True
  surfaces[floor_250] = True
  surfaces[floor_251] = True
  surfaces[floor_252] = True
  surfaces[floor_253] = True
  surfaces[floor_254] = True
  surfaces[floor_255] = True
  movable[couch_279] = True
  lieable[couch_279] = True
  surfaces[couch_279] = True
  sittable[couch_279] = True
  can_open[bookshelf_280] = True
  surfaces[bookshelf_280] = True
  containers[bookshelf_280] = True
  movable[table_281] = True
  surfaces[table_281] = True
  movable[desk_282] = True
  surfaces[desk_282] = True
  grabbable[chair_283] = True
  movable[chair_283] = True
  surfaces[chair_283] = True
  sittable[chair_283] = True
  can_open[dresser_284] = True
  containers[dresser_284] = True
  grabbable[hanger_285] = True
  movable[hanger_285] = True
  hangable[hanger_285] = True
  grabbable[hanger_287] = True
  movable[hanger_287] = True
  hangable[hanger_287] = True
  grabbable[hanger_289] = True
  movable[hanger_289] = True
  hangable[hanger_289] = True
  grabbable[hanger_291] = True
  movable[hanger_291] = True
  hangable[hanger_291] = True
  grabbable[hanger_293] = True
  movable[hanger_293] = True
  hangable[hanger_293] = True
  grabbable[hanger_295] = True
  movable[hanger_295] = True
  hangable[hanger_295] = True
  can_open[filing_cabinet_305] = True
  surfaces[filing_cabinet_305] = True
  containers[filing_cabinet_305] = True
  has_paper[drawing_307] = True
  cuttable[drawing_307] = True
  grabbable[drawing_307] = True
  movable[drawing_307] = True
  lookable[drawing_307] = True
  sittable[mat_308] = True
  grabbable[mat_308] = True
  movable[mat_308] = True
  lieable[mat_308] = True
  surfaces[mat_308] = True
  has_paper[drawing_309] = True
  cuttable[drawing_309] = True
  grabbable[drawing_309] = True
  movable[drawing_309] = True
  lookable[drawing_309] = True
  grabbable[pillow_310] = True
  movable[pillow_310] = True
  movable[curtain_311] = True
  can_open[curtain_311] = True
  cover_object[curtain_311] = True
  movable[curtain_312] = True
  can_open[curtain_312] = True
  cover_object[curtain_312] = True
  movable[curtain_313] = True
  can_open[curtain_313] = True
  cover_object[curtain_313] = True
  grabbable[toy_314] = True
  movable[toy_314] = True
  has_switch[television_315] = True
  lookable[television_315] = True
  has_plug[television_315] = True
  has_switch[light_316] = True
  has_plug[light_316] = True
  grabbable[mouse_318] = True
  movable[mouse_318] = True
  has_plug[mouse_318] = True
  movable[mousepad_319] = True
  surfaces[mousepad_319] = True
  lookable[computer_321] = True
  has_switch[computer_321] = True
  grabbable[keyboard_322] = True
  movable[keyboard_322] = True
  has_plug[keyboard_322] = True
  can_open[cupboard_1000] = True
  containers[cupboard_1000] = True
  grabbable[bowl_1001] = True
  movable[bowl_1001] = True
  recipient[bowl_1001] = True
  grabbable[food_oatmeal_1002] = True
  movable[food_oatmeal_1002] = True
  eatable[food_oatmeal_1002] = True
  pourable[milk_1003] = True
  grabbable[milk_1003] = True
  movable[milk_1003] = True
  drinkable[milk_1003] = True
  can_open[milk_1003] = True
  grabbable[ground_coffee_1004] = True
  movable[ground_coffee_1004] = True
  can_open[ground_coffee_1004] = True
  grabbable[cup_1005] = True
  movable[cup_1005] = True
  recipient[cup_1005] = True
  pourable[cup_1005] = True
  grabbable[juice_1006] = True
  movable[juice_1006] = True
  pourable[juice_1006] = True
  drinkable[juice_1006] = True
  grabbable[broom_2000] = True
  movable[broom_2000] = True
  grabbable[knife_2001] = True
  movable[knife_2001] = True
  grabbable[clothes_pants_2002] = True
  movable[clothes_pants_2002] = True
  clothes[clothes_pants_2002] = True
  hangable[clothes_pants_2002] = True
  pourable[blender_2003] = True
  grabbable[blender_2003] = True
  movable[blender_2003] = True
  recipient[blender_2003] = True
  has_switch[blender_2003] = True
  can_open[blender_2003] = True
  has_plug[blender_2003] = True
  grabbable[fork_2004] = True
  movable[fork_2004] = True
  grabbable[piano_bench_2005] = True
  movable[piano_bench_2005] = True
  surfaces[piano_bench_2005] = True
  sittable[piano_bench_2005] = True
  grabbable[pillow_2006] = True
  movable[pillow_2006] = True
  grabbable[shaving_cream_2007] = True
  movable[shaving_cream_2007] = True
  pourable[shaving_cream_2007] = True
  cream[shaving_cream_2007] = True
  grabbable[cup_2008] = True
  movable[cup_2008] = True
  recipient[cup_2008] = True
  pourable[cup_2008] = True
  grabbable[food_food_2009] = True
  movable[food_food_2009] = True
  eatable[food_food_2009] = True
  cuttable[food_food_2009] = True
  grabbable[clothes_skirt_2010] = True
  movable[clothes_skirt_2010] = True
  clothes[clothes_skirt_2010] = True
  hangable[clothes_skirt_2010] = True
  grabbable[towel_2011] = True
  movable[towel_2011] = True
  cover_object[towel_2011] = True
  grabbable[glue_2012] = True
  movable[glue_2012] = True
  cream[glue_2012] = True
  eatable[food_jam_2013] = True
  cream[food_jam_2013] = True
  grabbable[food_jam_2013] = True
  movable[food_jam_2013] = True
  can_open[food_jam_2013] = True
  has_paper[drawing_2014] = True
  cuttable[drawing_2014] = True
  grabbable[drawing_2014] = True
  movable[drawing_2014] = True
  lookable[drawing_2014] = True
  grabbable[food_food_2015] = True
  movable[food_food_2015] = True
  eatable[food_food_2015] = True
  cuttable[food_food_2015] = True
  grabbable[food_carrot_2016] = True
  movable[food_carrot_2016] = True
  eatable[food_carrot_2016] = True
  cuttable[food_carrot_2016] = True
  grabbable[comb_2017] = True
  movable[comb_2017] = True
  grabbable[stereo_2018] = True
  movable[stereo_2018] = True
  surfaces[stereo_2018] = True
  has_plug[stereo_2018] = True
  can_open[stereo_2018] = True
  has_switch[stereo_2018] = True
  grabbable[food_food_2019] = True
  movable[food_food_2019] = True
  eatable[food_food_2019] = True
  cuttable[food_food_2019] = True
  grabbable[band_aids_2020] = True
  movable[band_aids_2020] = True
  cuttable[band_aids_2020] = True
  grabbable[sheets_2021] = True
  movable[sheets_2021] = True
  cover_object[sheets_2021] = True
  containers[purse_2022] = True
  grabbable[purse_2022] = True
  movable[purse_2022] = True
  recipient[purse_2022] = True
  cover_object[purse_2022] = True
  can_open[purse_2022] = True
  grabbable[laundry_detergent_2023] = True
  movable[laundry_detergent_2023] = True
  pourable[laundry_detergent_2023] = True
  grabbable[food_food_2024] = True
  movable[food_food_2024] = True
  eatable[food_food_2024] = True
  cuttable[food_food_2024] = True
  grabbable[clothes_shirt_2025] = True
  movable[clothes_shirt_2025] = True
  clothes[clothes_shirt_2025] = True
  hangable[clothes_shirt_2025] = True
  grabbable[check_2026] = True
  movable[check_2026] = True
  readable[check_2026] = True
  has_paper[check_2026] = True
  grabbable[mouthwash_2027] = True
  movable[mouthwash_2027] = True
  pourable[mouthwash_2027] = True
  drinkable[mouthwash_2027] = True
  grabbable[video_game_controller_2028] = True
  movable[video_game_controller_2028] = True
  has_switch[video_game_controller_2028] = True
  has_plug[video_game_controller_2028] = True
  grabbable[form_2029] = True
  movable[form_2029] = True
  has_paper[form_2029] = True
  grabbable[needle_2030] = True
  movable[needle_2030] = True
  grabbable[button_2031] = True
  movable[button_2031] = True
  grabbable[wall_clock_2032] = True
  movable[wall_clock_2032] = True
  has_plug[wall_clock_2032] = True
  lookable[wall_clock_2032] = True
  has_switch[wall_clock_2032] = True
  grabbable[rag_2033] = True
  movable[rag_2033] = True
  recipient[rag_2033] = True
  cover_object[rag_2033] = True
  readable[novel_2034] = True
  cuttable[novel_2034] = True
  has_paper[novel_2034] = True
  grabbable[novel_2034] = True
  movable[novel_2034] = True
  can_open[novel_2034] = True
  grabbable[fork_2035] = True
  movable[fork_2035] = True
  grabbable[controller_2036] = True
  movable[controller_2036] = True
  has_plug[controller_2036] = True
  grabbable[centerpiece_2037] = True
  movable[centerpiece_2037] = True
  lookable[centerpiece_2037] = True
  cover_object[centerpiece_2037] = True
  grabbable[food_rice_2038] = True
  movable[food_rice_2038] = True
  pourable[food_rice_2038] = True
  eatable[food_rice_2038] = True
  grabbable[video_game_controller_2039] = True
  movable[video_game_controller_2039] = True
  has_switch[video_game_controller_2039] = True
  has_plug[video_game_controller_2039] = True
  grabbable[clothes_pants_2040] = True
  movable[clothes_pants_2040] = True
  clothes[clothes_pants_2040] = True
  hangable[clothes_pants_2040] = True
  grabbable[deck_of_cards_2041] = True
  movable[deck_of_cards_2041] = True
  has_paper[deck_of_cards_2041] = True
  readable[novel_2042] = True
  cuttable[novel_2042] = True
  has_paper[novel_2042] = True
  grabbable[novel_2042] = True
  movable[novel_2042] = True
  can_open[novel_2042] = True
  grabbable[juice_2043] = True
  movable[juice_2043] = True
  pourable[juice_2043] = True
  drinkable[juice_2043] = True
  grabbable[food_carrot_2044] = True
  movable[food_carrot_2044] = True
  eatable[food_carrot_2044] = True
  cuttable[food_carrot_2044] = True
  grabbable[check_2045] = True
  movable[check_2045] = True
  readable[check_2045] = True
  has_paper[check_2045] = True
  grabbable[ground_coffee_2046] = True
  movable[ground_coffee_2046] = True
  can_open[ground_coffee_2046] = True
  grabbable[piano_bench_2047] = True
  movable[piano_bench_2047] = True
  surfaces[piano_bench_2047] = True
  sittable[piano_bench_2047] = True
  pourable[blender_2048] = True
  grabbable[blender_2048] = True
  movable[blender_2048] = True
  recipient[blender_2048] = True
  has_switch[blender_2048] = True
  can_open[blender_2048] = True
  has_plug[blender_2048] = True
  grabbable[broom_2049] = True
  movable[broom_2049] = True
  grabbable[pencil_2050] = True
  movable[pencil_2050] = True
  grabbable[check_2051] = True
  movable[check_2051] = True
  readable[check_2051] = True
  has_paper[check_2051] = True
  grabbable[food_food_2052] = True
  movable[food_food_2052] = True
  eatable[food_food_2052] = True
  cuttable[food_food_2052] = True
  grabbable[oil_2053] = True
  movable[oil_2053] = True
  pourable[oil_2053] = True
  drinkable[oil_2053] = True
  grabbable[controller_2054] = True
  movable[controller_2054] = True
  has_plug[controller_2054] = True
  grabbable[food_food_2055] = True
  movable[food_food_2055] = True
  eatable[food_food_2055] = True
  cuttable[food_food_2055] = True
  grabbable[stamp_2056] = True
  movable[stamp_2056] = True
  grabbable[food_salt_2057] = True
  movable[food_salt_2057] = True
  pourable[food_salt_2057] = True
  eatable[food_salt_2057] = True
  grabbable[sheets_2058] = True
  movable[sheets_2058] = True
  cover_object[sheets_2058] = True
  grabbable[blow_dryer_2059] = True
  movable[blow_dryer_2059] = True
  has_switch[blow_dryer_2059] = True
  has_plug[blow_dryer_2059] = True
  grabbable[check_2060] = True
  movable[check_2060] = True
  readable[check_2060] = True
  has_paper[check_2060] = True
  containers[bag_2061] = True
  grabbable[bag_2061] = True
  movable[bag_2061] = True
  recipient[bag_2061] = True
  cover_object[bag_2061] = True
  can_open[bag_2061] = True
  grabbable[sheets_2062] = True
  movable[sheets_2062] = True
  cover_object[sheets_2062] = True
  grabbable[band_aids_2063] = True
  movable[band_aids_2063] = True
  cuttable[band_aids_2063] = True
  is_bathroom[bathroom_1]=True
  is_floor[floor_2]=True
  is_floor[floor_3]=True
  is_floor[floor_4]=True
  is_floor[floor_5]=True
  is_floor[floor_6]=True
  is_floor[floor_7]=True
  is_floor[floor_8]=True
  is_wall[wall_9]=True
  is_wall[wall_10]=True
  is_wall[wall_11]=True
  is_wall[wall_12]=True
  is_wall[wall_13]=True
  is_wall[wall_14]=True
  is_ceiling[ceiling_15]=True
  is_ceiling[ceiling_16]=True
  is_ceiling[ceiling_17]=True
  is_ceiling[ceiling_18]=True
  is_ceiling[ceiling_19]=True
  is_ceiling[ceiling_20]=True
  is_mat[mat_21]=True
  is_curtain[curtain_22]=True
  is_ceilinglamp[ceilinglamp_23]=True
  is_walllamp[walllamp_24]=True
  is_walllamp[walllamp_25]=True
  is_walllamp[walllamp_26]=True
  is_bathroom_counter[bathroom_counter_27]=True
  is_sink[sink_28]=True
  is_faucet[faucet_29]=True
  is_bathtub[bathtub_30]=True
  is_towel_rack[towel_rack_31]=True
  is_towel_rack[towel_rack_32]=True
  is_towel_rack[towel_rack_33]=True
  is_wallshelf[wallshelf_34]=True
  is_shower[shower_35]=True
  is_bathroom_cabinet[bathroom_cabinet_36]=True
  is_toilet[toilet_37]=True
  is_shelf[shelf_38]=True
  is_door[door_39]=True
  is_doorjamb[doorjamb_40]=True
  is_window[window_61]=True
  is_light[light_62]=True
  is_bedroom[bedroom_64]=True
  is_floor[floor_65]=True
  is_floor[floor_66]=True
  is_floor[floor_67]=True
  is_floor[floor_68]=True
  is_floor[floor_69]=True
  is_floor[floor_70]=True
  is_floor[floor_71]=True
  is_floor[floor_72]=True
  is_floor[floor_73]=True
  is_floor[floor_74]=True
  is_wall[wall_75]=True
  is_wall[wall_76]=True
  is_wall[wall_77]=True
  is_wall[wall_78]=True
  is_wall[wall_79]=True
  is_wall[wall_80]=True
  is_wall[wall_81]=True
  is_wall[wall_82]=True
  is_wall[wall_83]=True
  is_window[window_84]=True
  is_ceiling[ceiling_85]=True
  is_ceiling[ceiling_86]=True
  is_ceiling[ceiling_87]=True
  is_ceiling[ceiling_88]=True
  is_ceiling[ceiling_89]=True
  is_ceiling[ceiling_90]=True
  is_ceiling[ceiling_91]=True
  is_ceiling[ceiling_92]=True
  is_ceiling[ceiling_93]=True
  is_ceilinglamp[ceilinglamp_94]=True
  is_tablelamp[tablelamp_95]=True
  is_chair[chair_96]=True
  is_bookshelf[bookshelf_97]=True
  is_nightstand[nightstand_98]=True
  is_bed[bed_99]=True
  is_dresser[dresser_100]=True
  is_chair[chair_101]=True
  is_hanger[hanger_102]=True
  is_table[table_103]=True
  is_doorjamb[doorjamb_104]=True
  is_light[light_105]=True
  is_mat[mat_107]=True
  is_drawing[drawing_108]=True
  is_drawing[drawing_109]=True
  is_drawing[drawing_110]=True
  is_curtain[curtain_111]=True
  is_curtain[curtain_112]=True
  is_pillow[pillow_113]=True
  is_pillow[pillow_114]=True
  is_vase[vase_115]=True
  is_hanger[hanger_124]=True
  is_hanger[hanger_125]=True
  is_hanger[hanger_126]=True
  is_hanger[hanger_127]=True
  is_hanger[hanger_128]=True
  is_hanger[hanger_129]=True
  is_hanger[hanger_130]=True
  is_hanger[hanger_131]=True
  is_hanger[hanger_132]=True
  is_hanger[hanger_133]=True
  is_hanger[hanger_134]=True
  is_closetdrawer[closetdrawer_141]=True
  is_closetdrawer[closetdrawer_142]=True
  is_closetdrawer[closetdrawer_143]=True
  is_closetdrawer[closetdrawer_144]=True
  is_closetdrawer[closetdrawer_145]=True
  is_closetdrawer[closetdrawer_146]=True
  is_dining_room[dining_room_163]=True
  is_floor[floor_164]=True
  is_floor[floor_165]=True
  is_floor[floor_166]=True
  is_floor[floor_167]=True
  is_floor[floor_168]=True
  is_floor[floor_169]=True
  is_floor[floor_170]=True
  is_wall[wall_171]=True
  is_wall[wall_172]=True
  is_wall[wall_173]=True
  is_wall[wall_174]=True
  is_wall[wall_175]=True
  is_wall[wall_176]=True
  is_ceiling[ceiling_177]=True
  is_ceiling[ceiling_178]=True
  is_ceiling[ceiling_179]=True
  is_ceiling[ceiling_180]=True
  is_ceiling[ceiling_181]=True
  is_ceiling[ceiling_182]=True
  is_door[door_183]=True
  is_doorjamb[doorjamb_184]=True
  is_maindoor[maindoor_185]=True
  is_ceilinglamp[ceilinglamp_186]=True
  is_ceilinglamp[ceilinglamp_187]=True
  is_tvstand[tvstand_188]=True
  is_table[table_189]=True
  is_bench[bench_190]=True
  is_bench[bench_191]=True
  is_kitchen_counter[kitchen_counter_192]=True
  is_sink[sink_193]=True
  is_faucet[faucet_194]=True
  is_bookshelf[bookshelf_195]=True
  is_mat[mat_196]=True
  is_drawing[drawing_197]=True
  is_drawing[drawing_198]=True
  is_orchid[orchid_199]=True
  is_light[light_200]=True
  is_powersocket[powersocket_201]=True
  is_television[television_202]=True
  is_wall_clock[wall_clock_204]=True
  is_phone[phone_205]=True
  is_photoframe[photoframe_219]=True
  is_cutting_board[cutting_board_223]=True
  is_cutting_board[cutting_board_228]=True
  is_oven[oven_229]=True
  is_tray[tray_230]=True
  is_toaster[toaster_231]=True
  is_freezer[freezer_234]=True
  is_stovefan[stovefan_235]=True
  is_coffe_maker[coffe_maker_236]=True
  is_microwave[microwave_238]=True
  is_home_office[home_office_246]=True
  is_floor[floor_247]=True
  is_floor[floor_248]=True
  is_floor[floor_249]=True
  is_floor[floor_250]=True
  is_floor[floor_251]=True
  is_floor[floor_252]=True
  is_floor[floor_253]=True
  is_floor[floor_254]=True
  is_floor[floor_255]=True
  is_wall[wall_256]=True
  is_wall[wall_257]=True
  is_wall[wall_258]=True
  is_wall[wall_259]=True
  is_wall[wall_260]=True
  is_wall[wall_261]=True
  is_wall[wall_262]=True
  is_wall[wall_263]=True
  is_ceiling[ceiling_264]=True
  is_ceiling[ceiling_265]=True
  is_ceiling[ceiling_266]=True
  is_ceiling[ceiling_267]=True
  is_ceiling[ceiling_268]=True
  is_ceiling[ceiling_269]=True
  is_ceiling[ceiling_270]=True
  is_ceiling[ceiling_271]=True
  is_ceiling[ceiling_272]=True
  is_doorjamb[doorjamb_273]=True
  is_doorjamb[doorjamb_274]=True
  is_window[window_275]=True
  is_ceilinglamp[ceilinglamp_276]=True
  is_walllamp[walllamp_277]=True
  is_walllamp[walllamp_278]=True
  is_couch[couch_279]=True
  is_bookshelf[bookshelf_280]=True
  is_table[table_281]=True
  is_desk[desk_282]=True
  is_chair[chair_283]=True
  is_dresser[dresser_284]=True
  is_hanger[hanger_285]=True
  is_hanger[hanger_287]=True
  is_hanger[hanger_289]=True
  is_hanger[hanger_291]=True
  is_hanger[hanger_293]=True
  is_hanger[hanger_295]=True
  is_closetdrawer[closetdrawer_296]=True
  is_closetdrawer[closetdrawer_299]=True
  is_closetdrawer[closetdrawer_301]=True
  is_filing_cabinet[filing_cabinet_305]=True
  is_standingmirror[standingmirror_306]=True
  is_drawing[drawing_307]=True
  is_mat[mat_308]=True
  is_drawing[drawing_309]=True
  is_pillow[pillow_310]=True
  is_curtain[curtain_311]=True
  is_curtain[curtain_312]=True
  is_curtain[curtain_313]=True
  is_toy[toy_314]=True
  is_television[television_315]=True
  is_light[light_316]=True
  is_powersocket[powersocket_317]=True
  is_mouse[mouse_318]=True
  is_mousepad[mousepad_319]=True
  is_cpuscreen[cpuscreen_320]=True
  is_computer[computer_321]=True
  is_keyboard[keyboard_322]=True
  is_cupboard[cupboard_1000]=True
  is_bowl[bowl_1001]=True
  is_food_oatmeal[food_oatmeal_1002]=True
  is_milk[milk_1003]=True
  is_ground_coffee[ground_coffee_1004]=True
  is_cup[cup_1005]=True
  is_juice[juice_1006]=True
  is_broom[broom_2000]=True
  is_knife[knife_2001]=True
  is_clothes_pants[clothes_pants_2002]=True
  is_blender[blender_2003]=True
  is_fork[fork_2004]=True
  is_piano_bench[piano_bench_2005]=True
  is_pillow[pillow_2006]=True
  is_shaving_cream[shaving_cream_2007]=True
  is_cup[cup_2008]=True
  is_food_food[food_food_2009]=True
  is_clothes_skirt[clothes_skirt_2010]=True
  is_towel[towel_2011]=True
  is_glue[glue_2012]=True
  is_food_jam[food_jam_2013]=True
  is_drawing[drawing_2014]=True
  is_food_food[food_food_2015]=True
  is_food_carrot[food_carrot_2016]=True
  is_comb[comb_2017]=True
  is_stereo[stereo_2018]=True
  is_food_food[food_food_2019]=True
  is_band_aids[band_aids_2020]=True
  is_sheets[sheets_2021]=True
  is_purse[purse_2022]=True
  is_laundry_detergent[laundry_detergent_2023]=True
  is_food_food[food_food_2024]=True
  is_clothes_shirt[clothes_shirt_2025]=True
  is_check[check_2026]=True
  is_mouthwash[mouthwash_2027]=True
  is_video_game_controller[video_game_controller_2028]=True
  is_form[form_2029]=True
  is_needle[needle_2030]=True
  is_button[button_2031]=True
  is_wall_clock[wall_clock_2032]=True
  is_rag[rag_2033]=True
  is_novel[novel_2034]=True
  is_fork[fork_2035]=True
  is_controller[controller_2036]=True
  is_centerpiece[centerpiece_2037]=True
  is_food_rice[food_rice_2038]=True
  is_video_game_controller[video_game_controller_2039]=True
  is_clothes_pants[clothes_pants_2040]=True
  is_deck_of_cards[deck_of_cards_2041]=True
  is_novel[novel_2042]=True
  is_juice[juice_2043]=True
  is_food_carrot[food_carrot_2044]=True
  is_check[check_2045]=True
  is_ground_coffee[ground_coffee_2046]=True
  is_piano_bench[piano_bench_2047]=True
  is_blender[blender_2048]=True
  is_broom[broom_2049]=True
  is_pencil[pencil_2050]=True
  is_check[check_2051]=True
  is_food_food[food_food_2052]=True
  is_oil[oil_2053]=True
  is_controller[controller_2054]=True
  is_food_food[food_food_2055]=True
  is_stamp[stamp_2056]=True
  is_food_salt[food_salt_2057]=True
  is_sheets[sheets_2058]=True
  is_blow_dryer[blow_dryer_2059]=True
  is_check[check_2060]=True
  is_bag[bag_2061]=True
  is_sheets[sheets_2062]=True
  is_band_aids[band_aids_2063]=True
