Goal: Make a humburger
Additional information: You can make it by put raw tomato, cooked egg, raw onion, raw cheese, cooked bacon on a peace of raw bread, then put another peace of raw bread on the top.

behavior __goal__():
    body:
        bind bread1: item where:
            is_bread(bread1)
        bind bread2: item where:
            is_bread(bread2) and bread1 != bread2
        bind tomato: item where:
            is_tomato(tomato)
        bind egg: item where:
            is_egg(egg)
        bind onion: item where:
            is_onion(onion)
        bind cheese: item where:
            is_cheese(cheese)
        bind bacon: item where:
            is_bacon(bacon)
        achieve clean(tomato)
        achieve sliced(tomato)
        achieve clean(onion)
        achieve sliced(onion)
        achieve cooked(egg)
        achieve cooked(bacon)
        achieve on(tomato, bread1)
        achieve on(egg, tomato)
        achieve on(onion, egg)
        achieve on(cheese, onion)
        achieve on(bacon, cheese)
        achieve on(bread2, bacon)