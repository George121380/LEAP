domain "virtualhome"

typedef item: object
typedef character: object
typedef room: object

# Features without return type annotations are assumed to be returning boolean values.

#state
feature is_on(x: item)
feature is_off(x: item)
feature plugged(x: item)
feature unplugged(x: item)
feature open(x: item)
feature closed(x: item)
feature dirty(x: item)
feature clean(x: item)
feature sitting(x: character)
feature lying(x: character)

#add state
feature is_door(x: item)
feature is_explored(x: item)

#relationship
feature on(x: item, y: item)
feature inside(x: item, y: item)
feature between(x: item, y: item, z: item)
feature close_item(x: item, y: item)
feature close(x: character, y: item)
feature facing(x: item, y: item)
feature holds_rh(x: character, y: item)
feature holds_lh(x: character, y: item)

#Properties 
feature surfaces(x: item)
feature grabbable(x: item)
feature sittable(x: item)
feature lieable(x: item)
feature hangable(x: item)
feature drinkable(x: item)
feature eatable(x: item)
feature recipient(x: item)
feature cuttable(x: item)
feature pourable(x: item)
feature can_open(x: item)
feature has_switch(x: item)
feature readable(x: item)
feature lookable(x: item)
feature containers(x: item)
feature clothes(x: item)
feature person(x: item)
feature body_part(x: item)
feature cover_object(x: item)
feature has_plug(x: item)
feature has_paper(x: item)
feature movable(x: item)
feature cream(x: item)


object_constant char:character

#controllers
controller walk_executor(x: item)
controller switchoff_executor(x: item)
controller put_executor(x: item, y: item)
controller grab_executor(x: item)

#path problem is not considered

behavior walk(obj: item):
  goal: close(char, obj)
  body:
    walk_executor(obj)
  eff:
    close[char,obj] = True

behavior switch_off(obj: item):
  goal: is_off(obj)
  body:
    achieve close(char, obj)
    switchoff_executor(obj)
  eff:
    is_off[obj] = True
    is_on[obj] = False

def has_free_hand():
  symbol b = exists obj: item where: holds_rh(char, obj) or holds_lh(char, obj)
  symbol inverse_b = not b
  return inverse_b

behavior free_hand():
  goal: has_free_hand()
  body:
    if not has_free_hand():
      bind obj: item where: 
        surfaces(obj)
      bind inhand_obj: item where: 
        holds_rh(char, inhand_obj) or holds_lh(char, inhand_obj)
      put_executor(inhand_obj, obj)
  eff:
    if not has_free_hand():
      if holds_lh(char, inhand_obj):
        holds_lh[char, inhand_obj] = False
        on[inhand_obj,obj] = True
      else:
        holds_rh[char, inhand_obj] = False
        on[inhand_obj, obj] = True
      