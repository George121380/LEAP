 
def has_water_in_cup(cup:item):
    symbol has_water=exists o: item : is_water(o) and inside(o, cup)
    return has_water

behavior fill_cup_with_water(cup:item, faucet:item):
    body:
        achieve_once is_on(faucet)
        achieve has_water(cup)
        achieve_once is_off(faucet)

behavior __goal__():
    body:
        bind cup: item where:
            is_cup(cup) and id[cup]==2087
        bind faucet: item where:
            is_faucet(faucet) and id[faucet]==134
        fill_cup_with_water(cup, faucet)
