 
behavior wash_item(item:item):
    body:
        achieve_once clean(item)

behavior fill_pot_with_water(pot:item):
    body:
        achieve_once has_water(pot)

behavior cook_chicken(chicken:item, stove:item, pot:item):
    goal:
        achieve inside(chicken, pot)
    body:
        achieve_once is_on(stove)

behavior cut_ingredient(item:item, cutting_board:item):
    body:
        achieve_once on(item, cutting_board)
        achieve_once cut(item)

behavior __goal__():
    body:
        bind vegetable: item where:
            is_food_vegetable(vegetable)
        # Select vegetable item

        bind onion: item where:
            is_food_onion(onion)
        # Select onion item

        bind chicken: item where:
            is_food_chicken(chicken)
        # Select chicken item

        bind sink: item where:
            is_sink(sink)
        # Select a sink

        bind pot: item where:
            is_pot(pot)
        # Select a pot

        bind stove: item where:
            is_stove(stove)
        # Select a stove

        foreach item: item:
            if item == vegetable or item == onion or item == chicken:
                wash_item(item)
                # Wash all ingredients

        fill_pot_with_water(pot)
        cook_chicken(chicken, stove, pot)
        
        bind cutting_board: item where:
            is_cutting_board(cutting_board)
        # Select a cutting board

        foreach item: item:
            if item == vegetable or item == onion or item == chicken:
                cut_ingredient(item, cutting_board)
                # Cut all ingredients
