problem "virtualhome-problem"
domain "virtualhome.cdl"

#!pragma planner_is_goal_serializable=False
#!pragma planner_is_goal_ordered=True
#!pragma planner_always_commit_skeleton=True

objects:
  dining_room_1:item
  floor_2:item
  floor_3:item
  floor_4:item
  floor_5:item
  floor_6:item
  floor_7:item
  floor_8:item
  floor_9:item
  floor_10:item
  floor_11:item
  ceiling_12:item
  ceiling_13:item
  ceiling_14:item
  ceiling_15:item
  ceiling_16:item
  ceiling_17:item
  ceiling_18:item
  ceiling_19:item
  ceiling_20:item
  wall_21:item
  wall_22:item
  wall_23:item
  wall_24:item
  wall_25:item
  wall_26:item
  wall_27:item
  wall_28:item
  wall_29:item
  wall_30:item
  door_31:item
  doorjamb_32:item
  window_33:item
  ceilinglamp_34:item
  ceilinglamp_35:item
  walllamp_36:item
  chair_59:item
  chair_60:item
  chair_61:item
  chair_62:item
  table_63:item
  cupboard_64:item
  cupboard_65:item
  kitchen_counter_66:item
  sink_67:item
  faucet_68:item
  kitchen_counter_69:item
  kitchen_counter_70:item
  couch_71:item
  nightstand_72:item
  nightstand_73:item
  wallshelf_74:item
  wallshelf_75:item
  toaster_76:item
  stovefan_79:item
  freezer_80:item
  dishwasher_81:item
  oven_82:item
  tray_83:item
  coffe_maker_84:item
  microwave_86:item
  knifeblock_92:item
  pot_97:item
  pot_98:item
  photoframe_133:item
  mat_135:item
  orchid_136:item
  drawing_138:item
  drawing_139:item
  drawing_140:item
  drawing_141:item
  drawing_142:item
  curtain_143:item
  curtain_144:item
  curtain_145:item
  light_146:item
  powersocket_147:item
  phone_148:item
  bathroom_149:item
  wall_150:item
  wall_151:item
  wall_152:item
  wall_153:item
  ceiling_154:item
  ceiling_155:item
  ceiling_156:item
  ceiling_157:item
  floor_158:item
  floor_159:item
  floor_160:item
  floor_161:item
  floor_162:item
  walllamp_163:item
  ceilinglamp_164:item
  walllamp_165:item
  toilet_166:item
  shower_167:item
  bathroom_cabinet_168:item
  shower_169:item
  curtain_170:item
  bathroom_counter_171:item
  faucet_172:item
  sink_173:item
  mat_185:item
  drawing_186:item
  light_187:item
  bedroom_189:item
  bookshelf_190:item
  chair_191:item
  desk_192:item
  nightstand_193:item
  bed_194:item
  filing_cabinet_195:item
  light_196:item
  powersocket_197:item
  photoframe_204:item
  doorjamb_228:item
  door_229:item
  mat_230:item
  pillow_231:item
  pillow_232:item
  ceilinglamp_233:item
  floor_234:item
  floor_235:item
  floor_236:item
  floor_237:item
  floor_238:item
  ceiling_239:item
  ceiling_240:item
  ceiling_241:item
  ceiling_242:item
  wall_243:item
  wall_244:item
  wall_245:item
  wall_246:item
  home_office_248:item
  table_249:item
  bookshelf_250:item
  desk_251:item
  tvstand_252:item
  bookshelf_253:item
  chair_254:item
  nightstand_255:item
  couch_256:item
  couch_257:item
  dresser_258:item
  hanger_259:item
  hanger_260:item
  hanger_261:item
  hanger_262:item
  hanger_263:item
  hanger_264:item
  hanger_265:item
  closetdrawer_266:item
  closetdrawer_267:item
  closetdrawer_268:item
  closetdrawer_269:item
  closetdrawer_270:item
  closetdrawer_271:item
  closetdrawer_272:item
  computer_273:item
  cpuscreen_274:item
  keyboard_275:item
  mousepad_276:item
  mouse_277:item
  television_278:item
  powersocket_279:item
  light_280:item
  mat_281:item
  orchid_282:item
  drawing_283:item
  curtain_284:item
  curtain_285:item
  curtain_286:item
  pillow_287:item
  pillow_288:item
  pillow_289:item
  pillow_290:item
  photoframe_294:item
  ceilinglamp_310:item
  walllamp_311:item
  walllamp_312:item
  walllamp_313:item
  walllamp_314:item
  walllamp_315:item
  walllamp_316:item
  tablelamp_317:item
  wall_318:item
  wall_319:item
  wall_320:item
  wall_321:item
  wall_322:item
  wall_323:item
  wall_324:item
  wall_325:item
  ceiling_326:item
  ceiling_327:item
  ceiling_328:item
  ceiling_329:item
  ceiling_330:item
  ceiling_331:item
  ceiling_332:item
  ceiling_333:item
  ceiling_334:item
  floor_335:item
  floor_336:item
  floor_337:item
  floor_338:item
  floor_339:item
  floor_340:item
  floor_341:item
  floor_342:item
  floor_343:item
  floor_344:item
  doorjamb_345:item
  doorjamb_346:item
  door_347:item
  window_348:item
  kitchen_counter_1000:item
  cup_1001:item
  dishwasher_1002:item
  cup_1003:item
  plate_1004:item
  plate_1005:item
  dish_soap_1006:item
  dog_2000:item
  clothes_hat_2001:item
  check_2002:item
  check_2003:item
  clothes_scarf_2004:item
  oven_mitts_2005:item
  detergent_2006:item
  clothes_dress_2007:item
  food_food_2008:item
  needle_2009:item
  cup_2010:item
  cd_2011:item
  thread_2012:item
  shoe_rack_2013:item
  hanger_2014:item
  form_2015:item
  food_food_2016:item
  knife_2017:item
  food_carrot_2018:item
  napkin_2019:item
  soap_2020:item
  tray_2021:item
  food_peanut_butter_2022:item
  food_carrot_2023:item
  knife_2024:item
  cutting_board_2025:item
  juice_2026:item
  homework_2027:item
  clothes_hat_2028:item
  sponge_2029:item
  soap_2030:item
  food_food_2031:item
  sheets_2032:item
  food_food_2033:item
  toy_2034:item
  food_butter_2035:item
  pasta_2036:item
  soap_2037:item
  clothes_shirt_2038:item
  pencil_2039:item
  sponge_2040:item
  detergent_2041:item
  food_orange_2042:item
  sheets_2043:item
  tea_bag_2044:item
  food_food_2045:item
  bookmark_2046:item
  dvd_player_2047:item
  form_2048:item
  clothes_underwear_2049:item
  coffee_filter_2050:item
  newspaper_2051:item
  clothes_socks_2052:item
  bookmark_2053:item
  check_2054:item
  band_aids_2055:item
  detergent_2056:item
  keyboard_2057:item
  basket_for_clothes_2058:item
  toothbrush_holder_2059:item
  ground_coffee_2060:item
  toothbrush_holder_2061:item
  basket_for_clothes_2062:item
  after_shave_2063:item
  knife_2064:item
  food_food_2065:item
  shoes_2066:item
  wooden_spoon_2067:item
  char:character

init:
  clean[dining_room_1] = True
  is_room[dining_room_1]=True
  dirty[floor_2] = True
  clean[floor_3] = True
  clean[floor_4] = True
  dirty[floor_5] = True
  clean[floor_6] = True
  clean[floor_7] = True
  clean[floor_8] = True
  dirty[floor_9] = True
  dirty[floor_10] = True
  dirty[floor_11] = True
  dirty[ceiling_12] = True
  clean[ceiling_13] = True
  clean[ceiling_14] = True
  dirty[ceiling_15] = True
  dirty[ceiling_16] = True
  clean[ceiling_17] = True
  clean[ceiling_18] = True
  dirty[ceiling_19] = True
  clean[ceiling_20] = True
  clean[wall_21] = True
  clean[wall_22] = True
  clean[wall_23] = True
  clean[wall_24] = True
  dirty[wall_25] = True
  dirty[wall_26] = True
  clean[wall_27] = True
  clean[wall_28] = True
  dirty[wall_29] = True
  clean[wall_30] = True
  clean[door_31] = True
  open[door_31] = True
  clean[doorjamb_32] = True
  open[doorjamb_32] = True
  clean[window_33] = True
  open[window_33] = True
  clean[ceilinglamp_34] = True
  is_on[ceilinglamp_34] = True
  clean[ceilinglamp_35] = True
  is_on[ceilinglamp_35] = True
  clean[walllamp_36] = True
  is_on[walllamp_36] = True
  clean[chair_59] = True
  clean[chair_60] = True
  clean[chair_61] = True
  clean[chair_62] = True
  clean[table_63] = True
  clean[cupboard_64] = True
  open[cupboard_64] = True
  closed[cupboard_65] = True
  clean[cupboard_65] = True
  clean[kitchen_counter_66] = True
  open[kitchen_counter_66] = True
  clean[sink_67] = True
  clean[faucet_68] = True
  is_on[faucet_68] = True
  closed[kitchen_counter_69] = True
  clean[kitchen_counter_69] = True
  closed[kitchen_counter_70] = True
  clean[kitchen_counter_70] = True
  dirty[couch_71] = True
  clean[nightstand_72] = True
  open[nightstand_72] = True
  closed[nightstand_73] = True
  clean[nightstand_73] = True
  clean[wallshelf_74] = True
  clean[wallshelf_75] = True
  is_off[toaster_76] = True
  clean[toaster_76] = True
  plugged[toaster_76] = True
  clean[stovefan_79] = True
  clean[freezer_80] = True
  open[freezer_80] = True
  plugged[freezer_80] = True
  closed[dishwasher_81] = True
  clean[dishwasher_81] = True
  is_on[dishwasher_81] = True
  closed[oven_82] = True
  clean[oven_82] = True
  plugged[oven_82] = True
  is_off[oven_82] = True
  clean[tray_83] = True
  is_off[coffe_maker_84] = True
  clean[coffe_maker_84] = True
  open[coffe_maker_84] = True
  plugged[coffe_maker_84] = True
  closed[microwave_86] = True
  clean[microwave_86] = True
  plugged[microwave_86] = True
  is_off[microwave_86] = True
  clean[knifeblock_92] = True
  clean[pot_97] = True
  open[pot_97] = True
  closed[pot_98] = True
  dirty[pot_98] = True
  clean[photoframe_133] = True
  dirty[mat_135] = True
  clean[orchid_136] = True
  clean[drawing_138] = True
  clean[drawing_139] = True
  clean[drawing_140] = True
  clean[drawing_141] = True
  clean[drawing_142] = True
  closed[curtain_143] = True
  dirty[curtain_143] = True
  closed[curtain_144] = True
  clean[curtain_144] = True
  closed[curtain_145] = True
  dirty[curtain_145] = True
  clean[light_146] = True
  is_on[light_146] = True
  plugged[light_146] = True
  clean[powersocket_147] = True
  is_off[phone_148] = True
  clean[phone_148] = True
  plugged[phone_148] = True
  clean[bathroom_149] = True
  is_room[bathroom_149]=True
  clean[wall_150] = True
  clean[wall_151] = True
  clean[wall_152] = True
  dirty[wall_153] = True
  dirty[ceiling_154] = True
  clean[ceiling_155] = True
  dirty[ceiling_156] = True
  clean[ceiling_157] = True
  dirty[floor_158] = True
  clean[floor_159] = True
  clean[floor_160] = True
  clean[floor_161] = True
  dirty[floor_162] = True
  clean[walllamp_163] = True
  is_on[walllamp_163] = True
  clean[ceilinglamp_164] = True
  is_on[ceilinglamp_164] = True
  clean[walllamp_165] = True
  is_on[walllamp_165] = True
  is_off[toilet_166] = True
  clean[toilet_166] = True
  open[toilet_166] = True
  clean[shower_167] = True
  closed[bathroom_cabinet_168] = True
  clean[bathroom_cabinet_168] = True
  clean[shower_169] = True
  clean[curtain_170] = True
  open[curtain_170] = True
  clean[bathroom_counter_171] = True
  open[bathroom_counter_171] = True
  is_off[faucet_172] = True
  clean[faucet_172] = True
  clean[sink_173] = True
  clean[mat_185] = True
  clean[drawing_186] = True
  clean[light_187] = True
  is_on[light_187] = True
  plugged[light_187] = True
  clean[bedroom_189] = True
  is_room[bedroom_189]=True
  clean[bookshelf_190] = True
  open[bookshelf_190] = True
  clean[chair_191] = True
  clean[desk_192] = True
  clean[nightstand_193] = True
  open[nightstand_193] = True
  clean[bed_194] = True
  closed[filing_cabinet_195] = True
  clean[filing_cabinet_195] = True
  clean[light_196] = True
  is_on[light_196] = True
  plugged[light_196] = True
  clean[powersocket_197] = True
  clean[photoframe_204] = True
  clean[doorjamb_228] = True
  open[doorjamb_228] = True
  clean[door_229] = True
  open[door_229] = True
  dirty[mat_230] = True
  dirty[pillow_231] = True
  dirty[pillow_232] = True
  clean[ceilinglamp_233] = True
  is_on[ceilinglamp_233] = True
  clean[floor_234] = True
  dirty[floor_235] = True
  dirty[floor_236] = True
  dirty[floor_237] = True
  clean[floor_238] = True
  clean[ceiling_239] = True
  clean[ceiling_240] = True
  dirty[ceiling_241] = True
  dirty[ceiling_242] = True
  dirty[wall_243] = True
  dirty[wall_244] = True
  clean[wall_245] = True
  dirty[wall_246] = True
  clean[home_office_248] = True
  is_room[home_office_248]=True
  clean[table_249] = True
  closed[bookshelf_250] = True
  clean[bookshelf_250] = True
  clean[desk_251] = True
  clean[tvstand_252] = True
  closed[bookshelf_253] = True
  clean[bookshelf_253] = True
  clean[chair_254] = True
  clean[nightstand_255] = True
  open[nightstand_255] = True
  clean[couch_256] = True
  clean[couch_257] = True
  closed[dresser_258] = True
  clean[dresser_258] = True
  clean[hanger_259] = True
  clean[hanger_260] = True
  clean[hanger_261] = True
  clean[hanger_262] = True
  clean[hanger_263] = True
  clean[hanger_264] = True
  clean[hanger_265] = True
  clean[closetdrawer_266] = True
  clean[closetdrawer_267] = True
  clean[closetdrawer_268] = True
  clean[closetdrawer_269] = True
  clean[closetdrawer_270] = True
  clean[closetdrawer_271] = True
  clean[closetdrawer_272] = True
  is_off[computer_273] = True
  clean[computer_273] = True
  plugged[computer_273] = True
  clean[cpuscreen_274] = True
  clean[keyboard_275] = True
  unplugged[keyboard_275] = True
  dirty[mousepad_276] = True
  clean[mouse_277] = True
  plugged[mouse_277] = True
  is_off[television_278] = True
  clean[television_278] = True
  plugged[television_278] = True
  clean[powersocket_279] = True
  clean[light_280] = True
  is_on[light_280] = True
  plugged[light_280] = True
  clean[mat_281] = True
  clean[orchid_282] = True
  clean[drawing_283] = True
  closed[curtain_284] = True
  clean[curtain_284] = True
  clean[curtain_285] = True
  open[curtain_285] = True
  closed[curtain_286] = True
  clean[curtain_286] = True
  dirty[pillow_287] = True
  clean[pillow_288] = True
  clean[pillow_289] = True
  dirty[pillow_290] = True
  clean[photoframe_294] = True
  clean[ceilinglamp_310] = True
  is_on[ceilinglamp_310] = True
  clean[walllamp_311] = True
  is_on[walllamp_311] = True
  clean[walllamp_312] = True
  is_on[walllamp_312] = True
  clean[walllamp_313] = True
  is_on[walllamp_313] = True
  clean[walllamp_314] = True
  is_on[walllamp_314] = True
  clean[walllamp_315] = True
  is_on[walllamp_315] = True
  clean[walllamp_316] = True
  is_on[walllamp_316] = True
  clean[tablelamp_317] = True
  is_on[tablelamp_317] = True
  clean[wall_318] = True
  clean[wall_319] = True
  dirty[wall_320] = True
  clean[wall_321] = True
  clean[wall_322] = True
  dirty[wall_323] = True
  clean[wall_324] = True
  dirty[wall_325] = True
  dirty[ceiling_326] = True
  dirty[ceiling_327] = True
  dirty[ceiling_328] = True
  clean[ceiling_329] = True
  clean[ceiling_330] = True
  dirty[ceiling_331] = True
  dirty[ceiling_332] = True
  clean[ceiling_333] = True
  clean[ceiling_334] = True
  clean[floor_335] = True
  clean[floor_336] = True
  dirty[floor_337] = True
  dirty[floor_338] = True
  clean[floor_339] = True
  clean[floor_340] = True
  clean[floor_341] = True
  clean[floor_342] = True
  dirty[floor_343] = True
  dirty[floor_344] = True
  clean[doorjamb_345] = True
  open[doorjamb_345] = True
  clean[doorjamb_346] = True
  open[doorjamb_346] = True
  clean[door_347] = True
  open[door_347] = True
  clean[window_348] = True
  open[window_348] = True
  clean[kitchen_counter_1000] = True
  dirty[cup_1001] = True
  closed[dishwasher_1002] = True
  clean[dishwasher_1002] = True
  dirty[cup_1003] = True
  clean[plate_1004] = True
  clean[plate_1005] = True
  clean[dish_soap_1006] = True
  clean[dog_2000] = True
  clean[clothes_hat_2001] = True
  clean[check_2002] = True
  clean[check_2003] = True
  dirty[clothes_scarf_2004] = True
  clean[oven_mitts_2005] = True
  clean[detergent_2006] = True
  dirty[clothes_dress_2007] = True
  clean[food_food_2008] = True
  clean[needle_2009] = True
  dirty[cup_2010] = True
  clean[cd_2011] = True
  clean[thread_2012] = True
  clean[shoe_rack_2013] = True
  clean[hanger_2014] = True
  clean[form_2015] = True
  clean[food_food_2016] = True
  clean[knife_2017] = True
  dirty[food_carrot_2018] = True
  dirty[napkin_2019] = True
  clean[soap_2020] = True
  clean[tray_2021] = True
  clean[food_peanut_butter_2022] = True
  dirty[food_carrot_2023] = True
  clean[knife_2024] = True
  clean[cutting_board_2025] = True
  clean[juice_2026] = True
  clean[homework_2027] = True
  clean[clothes_hat_2028] = True
  dirty[sponge_2029] = True
  clean[soap_2030] = True
  clean[food_food_2031] = True
  clean[sheets_2032] = True
  dirty[food_food_2033] = True
  dirty[toy_2034] = True
  clean[food_butter_2035] = True
  clean[pasta_2036] = True
  clean[soap_2037] = True
  clean[clothes_shirt_2038] = True
  clean[pencil_2039] = True
  clean[sponge_2040] = True
  clean[detergent_2041] = True
  clean[food_orange_2042] = True
  dirty[sheets_2043] = True
  clean[tea_bag_2044] = True
  dirty[food_food_2045] = True
  clean[bookmark_2046] = True
  closed[dvd_player_2047] = True
  clean[dvd_player_2047] = True
  unplugged[dvd_player_2047] = True
  clean[form_2048] = True
  clean[clothes_underwear_2049] = True
  dirty[coffee_filter_2050] = True
  clean[newspaper_2051] = True
  open[newspaper_2051] = True
  clean[clothes_socks_2052] = True
  clean[bookmark_2053] = True
  clean[check_2054] = True
  clean[band_aids_2055] = True
  clean[detergent_2056] = True
  clean[keyboard_2057] = True
  plugged[keyboard_2057] = True
  clean[basket_for_clothes_2058] = True
  open[basket_for_clothes_2058] = True
  clean[toothbrush_holder_2059] = True
  clean[ground_coffee_2060] = True
  open[ground_coffee_2060] = True
  clean[toothbrush_holder_2061] = True
  clean[basket_for_clothes_2062] = True
  open[basket_for_clothes_2062] = True
  clean[after_shave_2063] = True
  open[after_shave_2063] = True
  clean[knife_2064] = True
  dirty[food_food_2065] = True
  clean[shoes_2066] = True
  clean[wooden_spoon_2067] = True
  close_item[food_carrot_2023,freezer_80]=True
  close_item[clothes_shirt_2038,couch_256]=True
  close_item[clothes_hat_2028,couch_71]=True
  close_item[sheets_2043,dresser_258]=True
  inside[freezer_80,dining_room_1]=True
  inside[detergent_2041,filing_cabinet_195]=True
  inside[detergent_2041,bedroom_189]=True
  inside[pillow_290,home_office_248]=True
  inside[pillow_290,couch_257]=True
  inside[ceiling_157,bathroom_149]=True
  close_item[computer_273,wall_322]=True
  close_item[computer_273,floor_344]=True
  close_item[computer_273,wall_325]=True
  close_item[computer_273,cpuscreen_274]=True
  close_item[computer_273,keyboard_275]=True
  close_item[computer_273,floor_339]=True
  close_item[computer_273,mousepad_276]=True
  close_item[computer_273,mouse_277]=True
  close_item[computer_273,floor_338]=True
  close_item[computer_273,walllamp_312]=True
  close_item[computer_273,desk_251]=True
  close_item[computer_273,chair_254]=True
  close_item[computer_273,wall_319]=True
  facing_item[floor_335,drawing_283]=True
  close_item[photoframe_294,wall_320]=True
  close_item[photoframe_294,wall_323]=True
  close_item[photoframe_294,ceiling_326]=True
  close_item[photoframe_294,floor_335]=True
  close_item[photoframe_294,floor_336]=True
  close_item[photoframe_294,wall_246]=True
  close_item[photoframe_294,bookshelf_253]=True
  inside[oven_mitts_2005,filing_cabinet_195]=True
  inside[oven_mitts_2005,bedroom_189]=True
  inside[cupboard_64,dining_room_1]=True
  close_item[walllamp_313,wall_323]=True
  close_item[walllamp_313,ceiling_326]=True
  close_item[walllamp_313,floor_335]=True
  close_item[walllamp_313,floor_336]=True
  close_item[walllamp_313,drawing_283]=True
  close_item[walllamp_313,bookshelf_253]=True
  close_item[walllamp_313,wall_318]=True
  close_item[wall_319,wall_322]=True
  close_item[wall_319,wall_325]=True
  close_item[wall_319,ceiling_329]=True
  close_item[wall_319,computer_273]=True
  close_item[wall_319,cpuscreen_274]=True
  close_item[wall_319,keyboard_275]=True
  close_item[wall_319,mousepad_276]=True
  close_item[wall_319,mouse_277]=True
  close_item[wall_319,floor_339]=True
  close_item[wall_319,walllamp_311]=True
  close_item[wall_319,walllamp_312]=True
  close_item[wall_319,doorjamb_346]=True
  close_item[wall_319,desk_251]=True
  close_item[ceiling_334,dresser_258]=True
  close_item[ceiling_334,hanger_259]=True
  close_item[ceiling_334,hanger_260]=True
  close_item[ceiling_334,hanger_261]=True
  close_item[ceiling_334,hanger_262]=True
  close_item[ceiling_334,hanger_263]=True
  close_item[ceiling_334,hanger_264]=True
  close_item[ceiling_334,hanger_265]=True
  close_item[ceiling_334,wall_325]=True
  close_item[ceiling_334,ceiling_329]=True
  close_item[ceiling_334,ceiling_333]=True
  close_item[ceiling_334,walllamp_312]=True
  close_item[ceiling_334,doorjamb_346]=True
  close_item[ceiling_334,walllamp_315]=True
  close_item[ceiling_334,curtain_284]=True
  close_item[ceiling_334,curtain_285]=True
  inside[form_2015,bedroom_189]=True
  close_item[wall_22,floor_2]=True
  close_item[wall_22,floor_3]=True
  close_item[wall_22,photoframe_133]=True
  close_item[wall_22,floor_6]=True
  close_item[wall_22,floor_5]=True
  close_item[wall_22,mat_135]=True
  close_item[wall_22,drawing_138]=True
  close_item[wall_22,drawing_139]=True
  close_item[wall_22,drawing_140]=True
  close_item[wall_22,drawing_141]=True
  close_item[wall_22,drawing_142]=True
  close_item[wall_22,ceiling_14]=True
  close_item[wall_22,ceiling_16]=True
  close_item[wall_22,ceiling_17]=True
  close_item[wall_22,light_146]=True
  close_item[wall_22,powersocket_147]=True
  close_item[wall_22,wall_23]=True
  close_item[wall_22,wall_153]=True
  close_item[wall_22,wall_28]=True
  close_item[wall_22,ceiling_156]=True
  close_item[wall_22,door_31]=True
  close_item[wall_22,doorjamb_32]=True
  close_item[wall_22,floor_161]=True
  close_item[wall_22,ceilinglamp_34]=True
  close_item[wall_22,toilet_166]=True
  close_item[wall_22,shower_167]=True
  close_item[wall_22,shower_169]=True
  close_item[wall_22,chair_59]=True
  close_item[wall_22,couch_71]=True
  close_item[wall_22,nightstand_73]=True
  close_item[wall_22,freezer_80]=True
  inside[wall_28,dining_room_1]=True
  inside[wall_325,home_office_248]=True
  close_item[wall_27,window_33]=True
  close_item[wall_27,floor_7]=True
  close_item[wall_27,wallshelf_74]=True
  close_item[wall_27,wallshelf_75]=True
  close_item[wall_27,curtain_143]=True
  close_item[wall_27,curtain_144]=True
  close_item[wall_27,curtain_145]=True
  close_item[wall_27,ceiling_18]=True
  close_item[wall_27,wall_29]=True
  close_item[wall_27,wall_30]=True
  inside[doorjamb_345,home_office_248]=True
  facing_item[floor_6,drawing_139]=True
  facing_item[floor_6,drawing_140]=True
  facing_item[floor_6,drawing_141]=True
  facing_item[floor_6,drawing_142]=True
  inside[computer_273,home_office_248]=True
  close_item[kitchen_counter_70,cupboard_64]=True
  close_item[kitchen_counter_70,soap_2020]=True
  close_item[kitchen_counter_70,kitchen_counter_69]=True
  close_item[kitchen_counter_70,floor_10]=True
  close_item[kitchen_counter_70,soap_2030]=True
  close_item[kitchen_counter_70,dishwasher_81]=True
  close_item[kitchen_counter_70,wooden_spoon_2067]=True
  close_item[kitchen_counter_70,coffe_maker_84]=True
  close_item[kitchen_counter_70,wall_25]=True
  close_item[kitchen_counter_70,wall_29]=True
  close_item[wallshelf_75,window_33]=True
  close_item[wallshelf_75,doorjamb_228]=True
  close_item[wallshelf_75,door_229]=True
  close_item[wallshelf_75,floor_8]=True
  close_item[wallshelf_75,wallshelf_74]=True
  close_item[wallshelf_75,curtain_143]=True
  close_item[wallshelf_75,curtain_144]=True
  close_item[wallshelf_75,ceiling_20]=True
  close_item[wallshelf_75,wall_27]=True
  close_item[wallshelf_75,wall_30]=True
  facing_item[pillow_288,drawing_283]=True
  facing_item[pillow_288,television_278]=True
  inside[nightstand_73,dining_room_1]=True
  inside[food_food_2008,home_office_248]=True
  inside[couch_257,home_office_248]=True
  inside[tea_bag_2044,cupboard_65]=True
  inside[tea_bag_2044,dining_room_1]=True
  on[freezer_80,floor_6]=True
  facing_item[photoframe_294,drawing_283]=True
  close_item[floor_337,wall_320]=True
  close_item[floor_337,couch_256]=True
  close_item[floor_337,wall_322]=True
  close_item[floor_337,filing_cabinet_195]=True
  close_item[floor_337,light_196]=True
  close_item[floor_337,wall_323]=True
  close_item[floor_337,mat_281]=True
  close_item[floor_337,floor_237]=True
  close_item[floor_337,floor_335]=True
  close_item[floor_337,floor_336]=True
  close_item[floor_337,floor_338]=True
  close_item[floor_337,floor_340]=True
  close_item[floor_337,wall_246]=True
  close_item[floor_337,powersocket_279]=True
  close_item[floor_337,light_280]=True
  close_item[floor_337,doorjamb_345]=True
  close_item[floor_337,bookshelf_250]=True
  close_item[floor_337,door_347]=True
  close_item[floor_337,bookshelf_253]=True
  close_item[floor_337,chair_254]=True
  close_item[wall_23,door_229]=True
  close_item[wall_23,doorjamb_228]=True
  close_item[wall_23,floor_5]=True
  close_item[wall_23,powersocket_197]=True
  close_item[wall_23,couch_71]=True
  close_item[wall_23,orchid_136]=True
  close_item[wall_23,nightstand_72]=True
  close_item[wall_23,drawing_138]=True
  close_item[wall_23,drawing_139]=True
  close_item[wall_23,drawing_140]=True
  close_item[wall_23,drawing_141]=True
  close_item[wall_23,drawing_142]=True
  close_item[wall_23,nightstand_73]=True
  close_item[wall_23,ceiling_16]=True
  close_item[wall_23,wall_243]=True
  close_item[wall_23,wall_22]=True
  close_item[wall_23,wall_30]=True
  inside[wall_21,dining_room_1]=True
  inside[wall_318,home_office_248]=True
  facing_item[faucet_172,drawing_186]=True
  on[toilet_166,floor_161]=True
  close_item[cupboard_65,ceiling_12]=True
  close_item[cupboard_65,ceiling_13]=True
  close_item[cupboard_65,phone_148]=True
  close_item[cupboard_65,wall_21]=True
  close_item[cupboard_65,wall_24]=True
  close_item[cupboard_65,wall_26]=True
  close_item[cupboard_65,walllamp_36]=True
  close_item[cupboard_65,kitchen_counter_66]=True
  close_item[cupboard_65,sink_67]=True
  close_item[cupboard_65,faucet_68]=True
  close_item[cupboard_65,toaster_76]=True
  close_item[cupboard_65,stovefan_79]=True
  close_item[cupboard_65,oven_82]=True
  close_item[cupboard_65,tray_83]=True
  close_item[cupboard_65,microwave_86]=True
  close_item[cupboard_65,knifeblock_92]=True
  close_item[cupboard_65,food_food_2016]=True
  close_item[cupboard_65,pot_97]=True
  close_item[cupboard_65,pot_98]=True
  close_item[cupboard_65,food_peanut_butter_2022]=True
  close_item[cupboard_65,knife_2024]=True
  close_item[cupboard_65,tea_bag_2044]=True
  inside[closetdrawer_266,home_office_248]=True
  inside[closetdrawer_266,dresser_258]=True
  on[tvstand_252,floor_343]=True
  inside[knifeblock_92,dining_room_1]=True
  close_item[wall_152,floor_161]=True
  close_item[wall_152,floor_162]=True
  close_item[wall_152,wall_153]=True
  close_item[wall_152,ceilinglamp_164]=True
  close_item[wall_152,walllamp_165]=True
  close_item[wall_152,ceiling_154]=True
  close_item[wall_152,bathroom_cabinet_168]=True
  close_item[wall_152,curtain_170]=True
  close_item[wall_152,bathroom_counter_171]=True
  close_item[wall_152,faucet_172]=True
  close_item[wall_152,sink_173]=True
  close_item[wall_152,wall_151]=True
  close_item[wall_152,mat_185]=True
  close_item[wall_152,drawing_186]=True
  close_item[wall_152,ceiling_156]=True
  close_item[wall_152,ceiling_157]=True
  close_item[wall_152,floor_158]=True
  close_item[wall_152,floor_159]=True
  inside[homework_2027,filing_cabinet_195]=True
  inside[homework_2027,bedroom_189]=True
  facing_item[wall_323,drawing_283]=True
  close_item[curtain_285,wall_321]=True
  close_item[curtain_285,dresser_258]=True
  close_item[curtain_285,hanger_259]=True
  close_item[curtain_285,hanger_260]=True
  close_item[curtain_285,wall_325]=True
  close_item[curtain_285,closetdrawer_267]=True
  close_item[curtain_285,closetdrawer_268]=True
  close_item[curtain_285,ceiling_333]=True
  close_item[curtain_285,ceiling_334]=True
  close_item[curtain_285,closetdrawer_271]=True
  close_item[curtain_285,tvstand_252]=True
  close_item[curtain_285,floor_343]=True
  close_item[curtain_285,television_278]=True
  close_item[curtain_285,window_348]=True
  close_item[curtain_285,walllamp_315]=True
  close_item[curtain_285,curtain_284]=True
  close_item[curtain_285,curtain_286]=True
  inside[toaster_76,dining_room_1]=True
  facing_item[door_347,computer_273]=True
  facing_item[door_347,drawing_283]=True
  close_item[walllamp_316,wall_321]=True
  close_item[walllamp_316,pillow_290]=True
  close_item[walllamp_316,couch_257]=True
  close_item[walllamp_316,wall_324]=True
  close_item[walllamp_316,ceiling_332]=True
  close_item[walllamp_316,ceiling_333]=True
  close_item[walllamp_316,floor_342]=True
  close_item[walllamp_316,table_249]=True
  close_item[walllamp_316,window_348]=True
  close_item[walllamp_316,curtain_286]=True
  inside[cd_2011,filing_cabinet_195]=True
  inside[cd_2011,bedroom_189]=True
  inside[floor_4,dining_room_1]=True
  inside[clothes_socks_2052,filing_cabinet_195]=True
  inside[clothes_socks_2052,bedroom_189]=True
  inside[wall_24,dining_room_1]=True
  inside[wall_321,home_office_248]=True
  facing_item[floor_337,computer_273]=True
  facing_item[floor_337,drawing_283]=True
  on[mat_185,floor_162]=True
  inside[wall_244,bedroom_189]=True
  inside[curtain_285,home_office_248]=True
  inside[curtain_285,curtain_284]=True
  close_item[chair_61,ceilinglamp_34]=True
  close_item[chair_61,floor_2]=True
  close_item[chair_61,floor_4]=True
  close_item[chair_61,floor_3]=True
  close_item[chair_61,floor_7]=True
  close_item[chair_61,floor_9]=True
  close_item[chair_61,floor_11]=True
  close_item[chair_61,wall_21]=True
  close_item[chair_61,chair_59]=True
  close_item[chair_61,chair_60]=True
  close_item[chair_61,chair_62]=True
  close_item[chair_61,table_63]=True
  close_item[kitchen_counter_66,cupboard_65]=True
  close_item[kitchen_counter_66,pot_98]=True
  close_item[kitchen_counter_66,sink_67]=True
  close_item[kitchen_counter_66,faucet_68]=True
  close_item[kitchen_counter_66,walllamp_36]=True
  close_item[kitchen_counter_66,pot_97]=True
  close_item[kitchen_counter_66,coffee_filter_2050]=True
  close_item[kitchen_counter_66,floor_9]=True
  close_item[kitchen_counter_66,floor_11]=True
  close_item[kitchen_counter_66,toaster_76]=True
  close_item[kitchen_counter_66,stovefan_79]=True
  close_item[kitchen_counter_66,oven_82]=True
  close_item[kitchen_counter_66,tray_83]=True
  close_item[kitchen_counter_66,phone_148]=True
  close_item[kitchen_counter_66,wall_21]=True
  close_item[kitchen_counter_66,microwave_86]=True
  close_item[kitchen_counter_66,wall_24]=True
  close_item[kitchen_counter_66,wall_26]=True
  close_item[kitchen_counter_66,knifeblock_92]=True
  close_item[walllamp_165,floor_162]=True
  close_item[walllamp_165,bathroom_cabinet_168]=True
  close_item[walllamp_165,bathroom_counter_171]=True
  close_item[walllamp_165,wall_152]=True
  close_item[walllamp_165,drawing_186]=True
  close_item[walllamp_165,ceiling_157]=True
  inside[desk_192,bedroom_189]=True
  inside[soap_2020,dining_room_1]=True
  inside[closetdrawer_269,home_office_248]=True
  inside[closetdrawer_269,dresser_258]=True
  inside[window_33,dining_room_1]=True
  on[cup_1003,kitchen_counter_1000]=True
  on[faucet_68,kitchen_counter_66]=True
  inside[bookshelf_253,home_office_248]=True
  close_item[floor_3,doorjamb_32]=True
  close_item[floor_3,floor_160]=True
  close_item[floor_3,floor_2]=True
  close_item[floor_3,floor_4]=True
  close_item[floor_3,toilet_166]=True
  close_item[floor_3,mat_135]=True
  close_item[floor_3,floor_6]=True
  close_item[floor_3,floor_9]=True
  close_item[floor_3,chair_59]=True
  close_item[floor_3,shower_167]=True
  close_item[floor_3,freezer_80]=True
  close_item[floor_3,light_146]=True
  close_item[floor_3,powersocket_147]=True
  close_item[floor_3,wall_21]=True
  close_item[floor_3,wall_22]=True
  close_item[floor_3,wall_150]=True
  close_item[floor_3,light_187]=True
  close_item[floor_3,wall_28]=True
  close_item[floor_3,chair_61]=True
  close_item[floor_3,door_31]=True
  facing_item[orchid_136,drawing_140]=True
  facing_item[orchid_136,drawing_141]=True
  close_item[newspaper_2051,couch_257]=True
  close_item[floor_8,nightstand_193]=True
  close_item[floor_8,doorjamb_228]=True
  close_item[floor_8,powersocket_197]=True
  close_item[floor_8,door_229]=True
  close_item[floor_8,floor_7]=True
  close_item[floor_8,orchid_136]=True
  close_item[floor_8,nightstand_72]=True
  close_item[floor_8,floor_5]=True
  close_item[floor_8,wallshelf_75]=True
  close_item[floor_8,floor_235]=True
  close_item[floor_8,floor_234]=True
  close_item[floor_8,pillow_231]=True
  close_item[floor_8,wall_243]=True
  close_item[floor_8,chair_60]=True
  close_item[floor_8,wall_30]=True
  close_item[detergent_2056,filing_cabinet_195]=True
  inside[floor_7,dining_room_1]=True
  on[bookshelf_190,floor_234]=True
  on[bookshelf_190,floor_235]=True
  facing_item[floor_160,drawing_186]=True
  on[ceiling_20,wall_30]=True
  close_item[form_2015,bookshelf_190]=True
  close_item[soap_2030,kitchen_counter_70]=True
  close_item[soap_2020,kitchen_counter_70]=True
  inside[television_278,home_office_248]=True
  close_item[food_butter_2035,microwave_86]=True
  inside[band_aids_2055,bathroom_149]=True
  close_item[shower_167,floor_2]=True
  close_item[shower_167,floor_3]=True
  close_item[shower_167,photoframe_133]=True
  close_item[shower_167,floor_6]=True
  close_item[shower_167,mat_135]=True
  close_item[shower_167,ceiling_14]=True
  close_item[shower_167,ceiling_17]=True
  close_item[shower_167,light_146]=True
  close_item[shower_167,powersocket_147]=True
  close_item[shower_167,wall_150]=True
  close_item[shower_167,wall_22]=True
  close_item[shower_167,wall_153]=True
  close_item[shower_167,ceiling_155]=True
  close_item[shower_167,ceiling_156]=True
  close_item[shower_167,wall_28]=True
  close_item[shower_167,door_31]=True
  close_item[shower_167,doorjamb_32]=True
  close_item[shower_167,floor_161]=True
  close_item[shower_167,floor_160]=True
  close_item[shower_167,ceilinglamp_164]=True
  close_item[shower_167,toilet_166]=True
  close_item[shower_167,shower_169]=True
  close_item[shower_167,curtain_170]=True
  close_item[shower_167,light_187]=True
  close_item[shower_167,freezer_80]=True
  close_item[faucet_172,floor_162]=True
  close_item[faucet_172,bathroom_cabinet_168]=True
  close_item[faucet_172,bathroom_counter_171]=True
  close_item[faucet_172,sink_173]=True
  close_item[faucet_172,wall_151]=True
  close_item[faucet_172,wall_152]=True
  close_item[faucet_172,mat_185]=True
  close_item[faucet_172,ceiling_154]=True
  close_item[faucet_172,ceiling_157]=True
  close_item[faucet_172,floor_158]=True
  close_item[faucet_172,floor_159]=True
  close_item[light_187,doorjamb_32]=True
  close_item[light_187,floor_160]=True
  close_item[light_187,floor_2]=True
  close_item[light_187,floor_3]=True
  close_item[light_187,mat_135]=True
  close_item[light_187,shower_167]=True
  close_item[light_187,floor_9]=True
  close_item[light_187,ceiling_13]=True
  close_item[light_187,ceiling_14]=True
  close_item[light_187,light_146]=True
  close_item[light_187,phone_148]=True
  close_item[light_187,wall_21]=True
  close_item[light_187,wall_150]=True
  close_item[light_187,ceiling_155]=True
  close_item[light_187,wall_28]=True
  close_item[light_187,door_31]=True
  close_item[hanger_265,dresser_258]=True
  close_item[hanger_265,hanger_259]=True
  close_item[hanger_265,hanger_260]=True
  close_item[hanger_265,hanger_261]=True
  close_item[hanger_265,hanger_262]=True
  close_item[hanger_265,hanger_263]=True
  close_item[hanger_265,hanger_264]=True
  close_item[hanger_265,wall_325]=True
  close_item[hanger_265,closetdrawer_266]=True
  close_item[hanger_265,closetdrawer_267]=True
  close_item[hanger_265,closetdrawer_269]=True
  close_item[hanger_265,ceiling_334]=True
  close_item[hanger_265,closetdrawer_270]=True
  close_item[hanger_265,doorjamb_346]=True
  close_item[hanger_265,walllamp_315]=True
  inside[mat_185,bathroom_149]=True
  close_item[curtain_286,wall_321]=True
  close_item[curtain_286,wall_324]=True
  close_item[curtain_286,ceiling_332]=True
  close_item[curtain_286,ceiling_333]=True
  close_item[curtain_286,walllamp_316]=True
  close_item[curtain_286,window_348]=True
  close_item[curtain_286,table_249]=True
  close_item[curtain_286,orchid_282]=True
  close_item[curtain_286,curtain_284]=True
  close_item[curtain_286,curtain_285]=True
  close_item[curtain_286,floor_343]=True
  on[ceiling_13,wall_21]=True
  on[toothbrush_holder_2061,bathroom_counter_171]=True
  on[keyboard_275,desk_251]=True
  on[clothes_underwear_2049,couch_257]=True
  inside[form_2048,filing_cabinet_195]=True
  inside[form_2048,bedroom_189]=True
  facing_item[pillow_289,television_278]=True
  close_item[ceiling_14,doorjamb_32]=True
  close_item[ceiling_14,ceilinglamp_34]=True
  close_item[ceiling_14,shower_167]=True
  close_item[ceiling_14,ceiling_155]=True
  close_item[ceiling_14,ceiling_13]=True
  close_item[ceiling_14,ceiling_15]=True
  close_item[ceiling_14,freezer_80]=True
  close_item[ceiling_14,ceiling_17]=True
  close_item[ceiling_14,light_146]=True
  close_item[ceiling_14,phone_148]=True
  close_item[ceiling_14,wall_21]=True
  close_item[ceiling_14,wall_22]=True
  close_item[ceiling_14,wall_150]=True
  close_item[ceiling_14,light_187]=True
  close_item[ceiling_14,wall_28]=True
  on[pasta_2036,table_63]=True
  close_item[basket_for_clothes_2062,mat_281]=True
  facing_item[floor_159,drawing_186]=True
  inside[ceiling_240,bedroom_189]=True
  close_item[chair_62,ceilinglamp_35]=True
  close_item[chair_62,floor_4]=True
  close_item[chair_62,floor_7]=True
  close_item[chair_62,floor_10]=True
  close_item[chair_62,floor_11]=True
  close_item[chair_62,wall_29]=True
  close_item[chair_62,chair_59]=True
  close_item[chair_62,chair_60]=True
  close_item[chair_62,chair_61]=True
  close_item[chair_62,table_63]=True
  close_item[sink_67,cupboard_65]=True
  close_item[sink_67,kitchen_counter_66]=True
  close_item[sink_67,faucet_68]=True
  close_item[sink_67,floor_9]=True
  close_item[sink_67,juice_2026]=True
  close_item[sink_67,floor_11]=True
  close_item[sink_67,toaster_76]=True
  close_item[sink_67,after_shave_2063]=True
  close_item[sink_67,wall_21]=True
  close_item[sink_67,microwave_86]=True
  close_item[sink_67,wall_24]=True
  close_item[sink_67,wall_26]=True
  close_item[sink_67,knifeblock_92]=True
  on[sponge_2029,kitchen_counter_69]=True
  inside[bathroom_cabinet_168,bathroom_149]=True
  close_item[food_food_2033,plate_1005]=True
  on[knife_2017,kitchen_counter_1000]=True
  inside[photoframe_204,bedroom_189]=True
  inside[photoframe_204,bookshelf_190]=True
  close_item[closetdrawer_272,dresser_258]=True
  close_item[closetdrawer_272,wall_325]=True
  close_item[closetdrawer_272,closetdrawer_266]=True
  close_item[closetdrawer_272,closetdrawer_267]=True
  close_item[closetdrawer_272,closetdrawer_268]=True
  close_item[closetdrawer_272,closetdrawer_269]=True
  close_item[closetdrawer_272,closetdrawer_270]=True
  close_item[closetdrawer_272,closetdrawer_271]=True
  close_item[closetdrawer_272,floor_344]=True
  close_item[closetdrawer_272,doorjamb_346]=True
  close_item[closetdrawer_272,walllamp_315]=True
  facing_item[sink_173,drawing_186]=True
  inside[wall_152,bathroom_149]=True
  close_item[pillow_231,nightstand_193]=True
  close_item[pillow_231,bed_194]=True
  close_item[pillow_231,mat_230]=True
  close_item[pillow_231,pillow_232]=True
  close_item[pillow_231,floor_8]=True
  close_item[pillow_231,floor_234]=True
  close_item[pillow_231,floor_235]=True
  close_item[pillow_231,floor_238]=True
  close_item[pillow_231,wall_243]=True
  close_item[pillow_231,wall_244]=True
  close_item[pillow_231,wall_30]=True
  close_item[wall_246,powersocket_279]=True
  close_item[wall_246,light_280]=True
  close_item[wall_246,mat_281]=True
  close_item[wall_246,photoframe_294]=True
  close_item[wall_246,chair_191]=True
  close_item[wall_246,wall_320]=True
  close_item[wall_246,desk_192]=True
  close_item[wall_246,bed_194]=True
  close_item[wall_246,filing_cabinet_195]=True
  close_item[wall_246,light_196]=True
  close_item[wall_246,ceiling_327]=True
  close_item[wall_246,floor_337]=True
  close_item[wall_246,doorjamb_345]=True
  close_item[wall_246,door_347]=True
  close_item[wall_246,mat_230]=True
  close_item[wall_246,ceilinglamp_233]=True
  close_item[wall_246,floor_236]=True
  close_item[wall_246,floor_237]=True
  close_item[wall_246,floor_238]=True
  close_item[wall_246,ceiling_240]=True
  close_item[wall_246,ceiling_241]=True
  close_item[wall_246,ceiling_242]=True
  close_item[wall_246,wall_244]=True
  close_item[wall_246,wall_245]=True
  close_item[wall_246,bookshelf_250]=True
  close_item[wall_246,bookshelf_253]=True
  inside[dishwasher_1002,bedroom_189]=True
  close_item[bookshelf_250,desk_192]=True
  close_item[bookshelf_250,wall_320]=True
  close_item[bookshelf_250,wall_322]=True
  close_item[bookshelf_250,filing_cabinet_195]=True
  close_item[bookshelf_250,mat_281]=True
  close_item[bookshelf_250,ceiling_327]=True
  close_item[bookshelf_250,ceiling_328]=True
  close_item[bookshelf_250,floor_236]=True
  close_item[bookshelf_250,floor_237]=True
  close_item[bookshelf_250,ceiling_240]=True
  close_item[bookshelf_250,floor_337]=True
  close_item[bookshelf_250,floor_338]=True
  close_item[bookshelf_250,wall_245]=True
  close_item[bookshelf_250,wall_246]=True
  close_item[bookshelf_250,light_280]=True
  close_item[bookshelf_250,doorjamb_345]=True
  close_item[bookshelf_250,door_347]=True
  close_item[ceiling_329,wall_322]=True
  close_item[ceiling_329,wall_325]=True
  close_item[ceiling_329,ceiling_328]=True
  close_item[ceiling_329,ceiling_330]=True
  close_item[ceiling_329,ceiling_334]=True
  close_item[ceiling_329,cpuscreen_274]=True
  close_item[ceiling_329,ceilinglamp_310]=True
  close_item[ceiling_329,walllamp_311]=True
  close_item[ceiling_329,walllamp_312]=True
  close_item[ceiling_329,wall_319]=True
  inside[table_249,home_office_248]=True
  on[drawing_139,wall_23]=True
  close_item[ceiling_15,ceilinglamp_34]=True
  close_item[ceiling_15,ceilinglamp_35]=True
  close_item[ceiling_15,ceiling_12]=True
  close_item[ceiling_15,ceiling_14]=True
  close_item[ceiling_15,ceiling_16]=True
  close_item[ceiling_15,ceiling_18]=True
  close_item[after_shave_2063,sink_67]=True
  on[door_347,floor_237]=True
  on[nightstand_73,floor_6]=True
  close_item[toy_2034,mat_230]=True
  inside[floor_161,bathroom_149]=True
  close_item[mouse_277,wall_322]=True
  close_item[mouse_277,floor_344]=True
  close_item[mouse_277,wall_325]=True
  close_item[mouse_277,computer_273]=True
  close_item[mouse_277,cpuscreen_274]=True
  close_item[mouse_277,keyboard_275]=True
  close_item[mouse_277,mousepad_276]=True
  close_item[mouse_277,floor_339]=True
  close_item[mouse_277,walllamp_312]=True
  close_item[mouse_277,desk_251]=True
  close_item[mouse_277,chair_254]=True
  close_item[mouse_277,wall_319]=True
  close_item[drawing_283,wall_323]=True
  close_item[drawing_283,ceiling_326]=True
  close_item[drawing_283,ceiling_331]=True
  close_item[drawing_283,floor_335]=True
  close_item[drawing_283,floor_336]=True
  close_item[drawing_283,floor_341]=True
  close_item[drawing_283,walllamp_313]=True
  close_item[drawing_283,walllamp_314]=True
  close_item[drawing_283,tablelamp_317]=True
  close_item[drawing_283,wall_318]=True
  close_item[drawing_283,nightstand_255]=True
  inside[bathroom_counter_171,bathroom_149]=True
  on[wall_25,kitchen_counter_69]=True
  facing_item[tvstand_252,computer_273]=True
  facing_item[tvstand_252,television_278]=True
  facing_item[floor_8,drawing_139]=True
  facing_item[floor_8,drawing_140]=True
  facing_item[floor_8,drawing_141]=True
  facing_item[floor_8,drawing_142]=True
  close_item[ceiling_331,couch_256]=True
  close_item[ceiling_331,wall_323]=True
  close_item[ceiling_331,wall_324]=True
  close_item[ceiling_331,ceiling_326]=True
  close_item[ceiling_331,ceiling_330]=True
  close_item[ceiling_331,ceiling_332]=True
  close_item[ceiling_331,ceilinglamp_310]=True
  close_item[ceiling_331,walllamp_314]=True
  close_item[ceiling_331,drawing_283]=True
  close_item[ceiling_331,tablelamp_317]=True
  close_item[ceiling_331,wall_318]=True
  inside[mat_135,dining_room_1]=True
  facing_item[doorjamb_32,drawing_141]=True
  close_item[floor_336,couch_256]=True
  close_item[floor_336,wall_323]=True
  close_item[floor_336,light_196]=True
  close_item[floor_336,photoframe_294]=True
  close_item[floor_336,mat_281]=True
  close_item[floor_336,floor_335]=True
  close_item[floor_336,floor_337]=True
  close_item[floor_336,door_347]=True
  close_item[floor_336,floor_341]=True
  close_item[floor_336,powersocket_279]=True
  close_item[floor_336,walllamp_313]=True
  close_item[floor_336,drawing_283]=True
  close_item[floor_336,bookshelf_253]=True
  close_item[floor_336,nightstand_255]=True
  close_item[ceiling_13,cupboard_65]=True
  close_item[ceiling_13,ceilinglamp_34]=True
  close_item[ceiling_13,faucet_68]=True
  close_item[ceiling_13,walllamp_36]=True
  close_item[ceiling_13,toaster_76]=True
  close_item[ceiling_13,ceiling_12]=True
  close_item[ceiling_13,ceiling_14]=True
  close_item[ceiling_13,stovefan_79]=True
  close_item[ceiling_13,phone_148]=True
  close_item[ceiling_13,wall_21]=True
  close_item[ceiling_13,microwave_86]=True
  close_item[ceiling_13,wall_24]=True
  close_item[ceiling_13,light_187]=True
  close_item[ceiling_13,knifeblock_92]=True
  close_item[toothbrush_holder_2061,bathroom_counter_171]=True
  close_item[ceiling_18,window_33]=True
  close_item[ceiling_18,ceilinglamp_35]=True
  close_item[ceiling_18,wallshelf_74]=True
  close_item[ceiling_18,curtain_143]=True
  close_item[ceiling_18,curtain_144]=True
  close_item[ceiling_18,curtain_145]=True
  close_item[ceiling_18,ceiling_15]=True
  close_item[ceiling_18,ceiling_19]=True
  close_item[ceiling_18,ceiling_20]=True
  close_item[ceiling_18,wall_27]=True
  close_item[ceiling_18,wall_29]=True
  close_item[ceiling_18,wall_30]=True
  close_item[window_33,wallshelf_74]=True
  close_item[window_33,wallshelf_75]=True
  close_item[window_33,curtain_143]=True
  close_item[window_33,curtain_144]=True
  close_item[window_33,curtain_145]=True
  close_item[window_33,ceiling_18]=True
  close_item[window_33,wall_27]=True
  close_item[window_33,wall_29]=True
  close_item[window_33,wall_30]=True
  close_item[shoes_2066,dresser_258]=True
  inside[walllamp_313,home_office_248]=True
  close_item[cupboard_64,pot_97]=True
  close_item[cupboard_64,pot_98]=True
  close_item[cupboard_64,napkin_2019]=True
  close_item[cupboard_64,walllamp_36]=True
  close_item[cupboard_64,kitchen_counter_69]=True
  close_item[cupboard_64,kitchen_counter_70]=True
  close_item[cupboard_64,ceiling_12]=True
  close_item[cupboard_64,stovefan_79]=True
  close_item[cupboard_64,dishwasher_81]=True
  close_item[cupboard_64,oven_82]=True
  close_item[cupboard_64,ceiling_19]=True
  close_item[cupboard_64,coffe_maker_84]=True
  close_item[cupboard_64,tray_83]=True
  close_item[cupboard_64,food_food_2065]=True
  close_item[cupboard_64,wall_25]=True
  close_item[cupboard_64,wall_26]=True
  close_item[cupboard_64,wall_29]=True
  close_item[food_food_2045,plate_1004]=True
  close_item[powersocket_279,wall_320]=True
  close_item[powersocket_279,filing_cabinet_195]=True
  close_item[powersocket_279,light_196]=True
  close_item[powersocket_279,wall_323]=True
  close_item[powersocket_279,mat_281]=True
  close_item[powersocket_279,floor_237]=True
  close_item[powersocket_279,floor_335]=True
  close_item[powersocket_279,floor_336]=True
  close_item[powersocket_279,floor_337]=True
  close_item[powersocket_279,wall_246]=True
  close_item[powersocket_279,light_280]=True
  close_item[powersocket_279,doorjamb_345]=True
  close_item[powersocket_279,door_347]=True
  close_item[powersocket_279,bookshelf_253]=True
  close_item[curtain_284,wall_321]=True
  close_item[curtain_284,dresser_258]=True
  close_item[curtain_284,hanger_259]=True
  close_item[curtain_284,hanger_260]=True
  close_item[curtain_284,wall_325]=True
  close_item[curtain_284,closetdrawer_267]=True
  close_item[curtain_284,closetdrawer_268]=True
  close_item[curtain_284,ceiling_333]=True
  close_item[curtain_284,ceiling_334]=True
  close_item[curtain_284,closetdrawer_271]=True
  close_item[curtain_284,tvstand_252]=True
  close_item[curtain_284,television_278]=True
  close_item[curtain_284,floor_343]=True
  close_item[curtain_284,walllamp_315]=True
  close_item[curtain_284,window_348]=True
  close_item[curtain_284,curtain_285]=True
  close_item[curtain_284,curtain_286]=True
  on[pillow_288,couch_256]=True
  facing_item[wall_320,computer_273]=True
  facing_item[wall_320,drawing_283]=True
  facing_item[floor_161,drawing_186]=True
  inside[ceilinglamp_164,bathroom_149]=True
  inside[clothes_shirt_2038,home_office_248]=True
  facing_item[door_31,drawing_141]=True
  facing_item[door_31,drawing_142]=True
  inside[window_348,home_office_248]=True
  on[pot_97,oven_82]=True
  inside[ceiling_332,home_office_248]=True
  close_item[drawing_139,couch_71]=True
  close_item[drawing_139,drawing_138]=True
  close_item[drawing_139,drawing_140]=True
  close_item[drawing_139,drawing_141]=True
  close_item[drawing_139,drawing_142]=True
  close_item[drawing_139,ceiling_16]=True
  close_item[drawing_139,ceiling_17]=True
  close_item[drawing_139,wall_22]=True
  close_item[drawing_139,wall_23]=True
  close_item[floor_159,floor_160]=True
  close_item[floor_159,floor_162]=True
  close_item[floor_159,walllamp_163]=True
  close_item[floor_159,bathroom_counter_171]=True
  close_item[floor_159,faucet_172]=True
  close_item[floor_159,sink_173]=True
  close_item[floor_159,wall_150]=True
  close_item[floor_159,wall_151]=True
  close_item[floor_159,wall_152]=True
  close_item[floor_159,mat_185]=True
  close_item[floor_159,floor_158]=True
  close_item[ceilinglamp_164,shower_167]=True
  close_item[ceilinglamp_164,shower_169]=True
  close_item[ceilinglamp_164,curtain_170]=True
  close_item[ceilinglamp_164,wall_150]=True
  close_item[ceilinglamp_164,wall_151]=True
  close_item[ceilinglamp_164,wall_152]=True
  close_item[ceilinglamp_164,wall_153]=True
  close_item[ceilinglamp_164,ceiling_154]=True
  close_item[ceilinglamp_164,ceiling_155]=True
  close_item[ceilinglamp_164,ceiling_156]=True
  close_item[ceilinglamp_164,ceiling_157]=True
  inside[dvd_player_2047,home_office_248]=True
  inside[light_280,home_office_248]=True
  facing_item[floor_343,computer_273]=True
  facing_item[floor_343,television_278]=True
  facing_item[curtain_170,drawing_186]=True
  inside[kitchen_counter_70,dining_room_1]=True
  close_item[wall_322,computer_273]=True
  close_item[wall_322,cpuscreen_274]=True
  close_item[wall_322,keyboard_275]=True
  close_item[wall_322,mousepad_276]=True
  close_item[wall_322,mouse_277]=True
  close_item[wall_322,light_280]=True
  close_item[wall_322,mat_281]=True
  close_item[wall_322,ceilinglamp_310]=True
  close_item[wall_322,walllamp_311]=True
  close_item[wall_322,wall_319]=True
  close_item[wall_322,desk_192]=True
  close_item[wall_322,wall_320]=True
  close_item[wall_322,filing_cabinet_195]=True
  close_item[wall_322,ceiling_327]=True
  close_item[wall_322,ceiling_328]=True
  close_item[wall_322,ceiling_329]=True
  close_item[wall_322,floor_337]=True
  close_item[wall_322,floor_338]=True
  close_item[wall_322,floor_339]=True
  close_item[wall_322,doorjamb_345]=True
  close_item[wall_322,door_347]=True
  close_item[wall_322,floor_236]=True
  close_item[wall_322,ceiling_240]=True
  close_item[wall_322,wall_245]=True
  close_item[wall_322,bookshelf_250]=True
  close_item[wall_322,desk_251]=True
  close_item[wall_322,chair_254]=True
  inside[food_food_2031,dining_room_1]=True
  close_item[floor_343,pillow_288]=True
  close_item[floor_343,wall_321]=True
  close_item[floor_343,couch_256]=True
  close_item[floor_343,wall_324]=True
  close_item[floor_343,wall_325]=True
  close_item[floor_343,closetdrawer_267]=True
  close_item[floor_343,closetdrawer_268]=True
  close_item[floor_343,closetdrawer_271]=True
  close_item[floor_343,floor_340]=True
  close_item[floor_343,curtain_284]=True
  close_item[floor_343,television_278]=True
  close_item[floor_343,window_348]=True
  close_item[floor_343,floor_344]=True
  close_item[floor_343,table_249]=True
  close_item[floor_343,orchid_282]=True
  close_item[floor_343,floor_342]=True
  close_item[floor_343,tvstand_252]=True
  close_item[floor_343,curtain_285]=True
  close_item[floor_343,curtain_286]=True
  close_item[floor_343,pillow_287]=True
  on[plate_1004,kitchen_counter_1000]=True
  inside[floor_341,home_office_248]=True
  inside[pillow_289,home_office_248]=True
  close_item[cutting_board_2025,table_63]=True
  inside[stovefan_79,dining_room_1]=True
  close_item[hanger_264,dresser_258]=True
  close_item[hanger_264,hanger_259]=True
  close_item[hanger_264,hanger_260]=True
  close_item[hanger_264,hanger_261]=True
  close_item[hanger_264,hanger_262]=True
  close_item[hanger_264,hanger_263]=True
  close_item[hanger_264,wall_325]=True
  close_item[hanger_264,hanger_265]=True
  close_item[hanger_264,closetdrawer_266]=True
  close_item[hanger_264,closetdrawer_267]=True
  close_item[hanger_264,closetdrawer_269]=True
  close_item[hanger_264,ceiling_334]=True
  close_item[hanger_264,closetdrawer_270]=True
  close_item[hanger_264,doorjamb_346]=True
  inside[drawing_140,dining_room_1]=True
  inside[hanger_2014,home_office_248]=True
  inside[hanger_263,home_office_248]=True
  inside[hanger_263,dresser_258]=True
  on[mousepad_276,desk_251]=True
  close_item[floor_238,nightstand_193]=True
  close_item[floor_238,bed_194]=True
  close_item[floor_238,door_229]=True
  close_item[floor_238,mat_230]=True
  close_item[floor_238,pillow_231]=True
  close_item[floor_238,pillow_232]=True
  close_item[floor_238,floor_234]=True
  close_item[floor_238,floor_235]=True
  close_item[floor_238,floor_237]=True
  close_item[floor_238,wall_243]=True
  close_item[floor_238,wall_244]=True
  close_item[floor_238,wall_246]=True
  inside[toy_2034,bedroom_189]=True
  facing_item[television_278,computer_273]=True
  on[coffee_filter_2050,kitchen_counter_66]=True
  inside[table_63,dining_room_1]=True
  inside[floor_344,home_office_248]=True
  inside[floor_11,dining_room_1]=True
  facing_item[ceiling_156,drawing_186]=True
  inside[toothbrush_holder_2059,filing_cabinet_195]=True
  inside[toothbrush_holder_2059,bedroom_189]=True
  facing_item[bookshelf_253,drawing_283]=True
  on[closetdrawer_269,closetdrawer_270]=True
  inside[ceiling_328,home_office_248]=True
  facing_item[closetdrawer_271,computer_273]=True
  close_item[clothes_hat_2001,couch_71]=True
  close_item[tray_2021,couch_256]=True
  close_item[juice_2026,sink_67]=True
  inside[couch_256,home_office_248]=True
  close_item[sheets_2032,bed_194]=True
  inside[oven_82,dining_room_1]=True
  inside[sheets_2043,home_office_248]=True
  inside[sheets_2043,dresser_258]=True
  on[food_carrot_2018,plate_1004]=True
  facing_item[ceiling_331,drawing_283]=True
  facing_item[ceiling_331,television_278]=True
  inside[clothes_dress_2007,home_office_248]=True
  inside[kitchen_counter_66,dining_room_1]=True
  inside[ceiling_20,dining_room_1]=True
  close_item[wall_323,couch_256]=True
  close_item[wall_323,powersocket_279]=True
  close_item[wall_323,mat_281]=True
  close_item[wall_323,drawing_283]=True
  close_item[wall_323,pillow_288]=True
  close_item[wall_323,photoframe_294]=True
  close_item[wall_323,ceilinglamp_310]=True
  close_item[wall_323,walllamp_313]=True
  close_item[wall_323,walllamp_314]=True
  close_item[wall_323,tablelamp_317]=True
  close_item[wall_323,wall_318]=True
  close_item[wall_323,wall_320]=True
  close_item[wall_323,light_196]=True
  close_item[wall_323,ceiling_326]=True
  close_item[wall_323,ceiling_327]=True
  close_item[wall_323,ceiling_331]=True
  close_item[wall_323,floor_335]=True
  close_item[wall_323,floor_336]=True
  close_item[wall_323,floor_337]=True
  close_item[wall_323,floor_341]=True
  close_item[wall_323,doorjamb_345]=True
  close_item[wall_323,door_347]=True
  close_item[wall_323,bookshelf_253]=True
  close_item[wall_323,nightstand_255]=True
  close_item[ceiling_241,wall_320]=True
  close_item[ceiling_241,light_196]=True
  close_item[ceiling_241,ceiling_327]=True
  close_item[ceiling_241,ceilinglamp_233]=True
  close_item[ceiling_241,ceiling_240]=True
  close_item[ceiling_241,ceiling_242]=True
  close_item[ceiling_241,wall_244]=True
  close_item[ceiling_241,wall_245]=True
  close_item[ceiling_241,wall_246]=True
  close_item[ceiling_241,light_280]=True
  close_item[ceiling_241,doorjamb_345]=True
  close_item[ceiling_328,wall_322]=True
  close_item[ceiling_328,ceiling_327]=True
  close_item[ceiling_328,ceiling_329]=True
  close_item[ceiling_328,ceiling_240]=True
  close_item[ceiling_328,cpuscreen_274]=True
  close_item[ceiling_328,wall_245]=True
  close_item[ceiling_328,ceilinglamp_310]=True
  close_item[ceiling_328,walllamp_311]=True
  close_item[ceiling_328,bookshelf_250]=True
  on[drawing_140,wall_23]=True
  inside[clothes_hat_2001,dining_room_1]=True
  close_item[floor_5,floor_4]=True
  close_item[floor_5,powersocket_197]=True
  close_item[floor_5,floor_6]=True
  close_item[floor_5,couch_71]=True
  close_item[floor_5,nightstand_72]=True
  close_item[floor_5,orchid_136]=True
  close_item[floor_5,floor_8]=True
  close_item[floor_5,nightstand_73]=True
  close_item[floor_5,door_229]=True
  close_item[floor_5,wall_22]=True
  close_item[floor_5,wall_23]=True
  close_item[floor_5,chair_59]=True
  close_item[floor_5,chair_60]=True
  close_item[floor_5,wall_30]=True
  close_item[floor_5,table_63]=True
  close_item[bookmark_2053,desk_192]=True
  inside[wall_30,dining_room_1]=True
  inside[ceiling_327,home_office_248]=True
  close_item[floor_10,kitchen_counter_69]=True
  close_item[floor_10,kitchen_counter_70]=True
  close_item[floor_10,floor_7]=True
  close_item[floor_10,floor_11]=True
  close_item[floor_10,dishwasher_81]=True
  close_item[floor_10,coffe_maker_84]=True
  close_item[floor_10,wall_25]=True
  close_item[floor_10,wall_29]=True
  close_item[floor_10,chair_62]=True
  close_item[wall_25,cupboard_64]=True
  close_item[wall_25,pot_97]=True
  close_item[wall_25,pot_98]=True
  close_item[wall_25,walllamp_36]=True
  close_item[wall_25,kitchen_counter_69]=True
  close_item[wall_25,kitchen_counter_70]=True
  close_item[wall_25,floor_10]=True
  close_item[wall_25,ceiling_12]=True
  close_item[wall_25,stovefan_79]=True
  close_item[wall_25,dishwasher_81]=True
  close_item[wall_25,oven_82]=True
  close_item[wall_25,ceiling_19]=True
  close_item[wall_25,coffe_maker_84]=True
  close_item[wall_25,tray_83]=True
  close_item[wall_25,wall_26]=True
  close_item[wall_25,wall_29]=True
  facing_item[wall_321,television_278]=True
  close_item[basket_for_clothes_2058,dresser_258]=True
  on[newspaper_2051,couch_257]=True
  inside[floor_234,bedroom_189]=True
  close_item[soap_2037,sink_173]=True
  inside[walllamp_311,home_office_248]=True
  close_item[closetdrawer_271,wall_321]=True
  close_item[closetdrawer_271,dresser_258]=True
  close_item[closetdrawer_271,wall_325]=True
  close_item[closetdrawer_271,closetdrawer_266]=True
  close_item[closetdrawer_271,closetdrawer_267]=True
  close_item[closetdrawer_271,closetdrawer_268]=True
  close_item[closetdrawer_271,closetdrawer_269]=True
  close_item[closetdrawer_271,closetdrawer_270]=True
  close_item[closetdrawer_271,closetdrawer_272]=True
  close_item[closetdrawer_271,tvstand_252]=True
  close_item[closetdrawer_271,window_348]=True
  close_item[closetdrawer_271,television_278]=True
  close_item[closetdrawer_271,floor_343]=True
  close_item[closetdrawer_271,floor_344]=True
  close_item[closetdrawer_271,walllamp_315]=True
  close_item[closetdrawer_271,curtain_284]=True
  close_item[closetdrawer_271,curtain_285]=True
  inside[wallshelf_75,dining_room_1]=True
  close_item[mousepad_276,wall_322]=True
  close_item[mousepad_276,wall_325]=True
  close_item[mousepad_276,computer_273]=True
  close_item[mousepad_276,cpuscreen_274]=True
  close_item[mousepad_276,keyboard_275]=True
  close_item[mousepad_276,floor_339]=True
  close_item[mousepad_276,mouse_277]=True
  close_item[mousepad_276,walllamp_312]=True
  close_item[mousepad_276,desk_251]=True
  close_item[mousepad_276,chair_254]=True
  close_item[mousepad_276,wall_319]=True
  inside[cup_2010,home_office_248]=True
  inside[hanger_259,home_office_248]=True
  inside[hanger_259,dresser_258]=True
  facing_item[floor_340,computer_273]=True
  facing_item[floor_340,drawing_283]=True
  inside[chair_59,dining_room_1]=True
  inside[wall_243,bedroom_189]=True
  close_item[ceiling_12,cupboard_64]=True
  close_item[ceiling_12,pot_97]=True
  close_item[ceiling_12,pot_98]=True
  close_item[ceiling_12,cupboard_65]=True
  close_item[ceiling_12,walllamp_36]=True
  close_item[ceiling_12,ceilinglamp_34]=True
  close_item[ceiling_12,ceilinglamp_35]=True
  close_item[ceiling_12,toaster_76]=True
  close_item[ceiling_12,ceiling_13]=True
  close_item[ceiling_12,stovefan_79]=True
  close_item[ceiling_12,ceiling_15]=True
  close_item[ceiling_12,oven_82]=True
  close_item[ceiling_12,ceiling_19]=True
  close_item[ceiling_12,wall_21]=True
  close_item[ceiling_12,wall_24]=True
  close_item[ceiling_12,wall_25]=True
  close_item[ceiling_12,wall_26]=True
  close_item[ceiling_12,knifeblock_92]=True
  close_item[ceiling_12,wall_29]=True
  close_item[ground_coffee_2060,coffe_maker_84]=True
  inside[wall_23,dining_room_1]=True
  facing_item[curtain_144,drawing_139]=True
  facing_item[curtain_144,drawing_140]=True
  close_item[doorjamb_32,floor_160]=True
  close_item[doorjamb_32,floor_2]=True
  close_item[doorjamb_32,floor_3]=True
  close_item[doorjamb_32,toilet_166]=True
  close_item[doorjamb_32,mat_135]=True
  close_item[doorjamb_32,shower_167]=True
  close_item[doorjamb_32,ceiling_155]=True
  close_item[doorjamb_32,ceiling_14]=True
  close_item[doorjamb_32,freezer_80]=True
  close_item[doorjamb_32,light_146]=True
  close_item[doorjamb_32,powersocket_147]=True
  close_item[doorjamb_32,phone_148]=True
  close_item[doorjamb_32,wall_21]=True
  close_item[doorjamb_32,wall_150]=True
  close_item[doorjamb_32,wall_22]=True
  close_item[doorjamb_32,wall_153]=True
  close_item[doorjamb_32,light_187]=True
  close_item[doorjamb_32,wall_28]=True
  close_item[doorjamb_32,door_31]=True
  close_item[pencil_2039,table_249]=True
  inside[closetdrawer_268,home_office_248]=True
  inside[closetdrawer_268,dresser_258]=True
  close_item[kitchen_counter_69,cupboard_64]=True
  close_item[kitchen_counter_69,pot_97]=True
  close_item[kitchen_counter_69,pot_98]=True
  close_item[kitchen_counter_69,walllamp_36]=True
  close_item[kitchen_counter_69,kitchen_counter_70]=True
  close_item[kitchen_counter_69,floor_10]=True
  close_item[kitchen_counter_69,floor_11]=True
  close_item[kitchen_counter_69,sponge_2029]=True
  close_item[kitchen_counter_69,stovefan_79]=True
  close_item[kitchen_counter_69,food_food_2031]=True
  close_item[kitchen_counter_69,dishwasher_81]=True
  close_item[kitchen_counter_69,oven_82]=True
  close_item[kitchen_counter_69,tray_83]=True
  close_item[kitchen_counter_69,coffe_maker_84]=True
  close_item[kitchen_counter_69,wall_25]=True
  close_item[kitchen_counter_69,wall_26]=True
  close_item[kitchen_counter_69,wall_29]=True
  close_item[tea_bag_2044,cupboard_65]=True
  inside[sponge_2029,dining_room_1]=True
  inside[chair_191,bedroom_189]=True
  close_item[cpuscreen_274,wall_322]=True
  close_item[cpuscreen_274,ceiling_328]=True
  close_item[cpuscreen_274,ceiling_329]=True
  close_item[cpuscreen_274,computer_273]=True
  close_item[cpuscreen_274,floor_338]=True
  close_item[cpuscreen_274,keyboard_275]=True
  close_item[cpuscreen_274,mousepad_276]=True
  close_item[cpuscreen_274,mouse_277]=True
  close_item[cpuscreen_274,floor_339]=True
  close_item[cpuscreen_274,walllamp_311]=True
  close_item[cpuscreen_274,walllamp_312]=True
  close_item[cpuscreen_274,desk_251]=True
  close_item[cpuscreen_274,chair_254]=True
  close_item[cpuscreen_274,wall_319]=True
  close_item[pillow_289,couch_256]=True
  close_item[pillow_289,couch_257]=True
  close_item[pillow_289,pillow_290]=True
  close_item[pillow_289,wall_324]=True
  close_item[pillow_289,ceiling_332]=True
  close_item[pillow_289,floor_341]=True
  close_item[pillow_289,floor_342]=True
  close_item[pillow_289,tablelamp_317]=True
  close_item[pillow_289,wall_318]=True
  close_item[pillow_289,nightstand_255]=True
  close_item[ceilinglamp_310,couch_256]=True
  close_item[ceilinglamp_310,wall_322]=True
  close_item[ceilinglamp_310,wall_323]=True
  close_item[ceilinglamp_310,ceiling_326]=True
  close_item[ceilinglamp_310,ceiling_327]=True
  close_item[ceilinglamp_310,ceiling_328]=True
  close_item[ceilinglamp_310,ceiling_329]=True
  close_item[ceilinglamp_310,ceiling_330]=True
  close_item[ceilinglamp_310,ceiling_331]=True
  inside[check_2003,home_office_248]=True
  close_item[walllamp_314,couch_256]=True
  close_item[walllamp_314,couch_257]=True
  close_item[walllamp_314,wall_323]=True
  close_item[walllamp_314,ceiling_326]=True
  close_item[walllamp_314,ceiling_331]=True
  close_item[walllamp_314,floor_341]=True
  close_item[walllamp_314,drawing_283]=True
  close_item[walllamp_314,tablelamp_317]=True
  close_item[walllamp_314,wall_318]=True
  close_item[walllamp_314,nightstand_255]=True
  close_item[floor_335,couch_256]=True
  close_item[floor_335,wall_323]=True
  close_item[floor_335,light_196]=True
  close_item[floor_335,photoframe_294]=True
  close_item[floor_335,mat_281]=True
  close_item[floor_335,floor_336]=True
  close_item[floor_335,floor_337]=True
  close_item[floor_335,door_347]=True
  close_item[floor_335,floor_341]=True
  close_item[floor_335,powersocket_279]=True
  close_item[floor_335,walllamp_313]=True
  close_item[floor_335,drawing_283]=True
  close_item[floor_335,bookshelf_253]=True
  close_item[floor_335,nightstand_255]=True
  inside[floor_6,dining_room_1]=True
  inside[check_2054,filing_cabinet_195]=True
  inside[check_2054,bedroom_189]=True
  facing_item[curtain_143,drawing_139]=True
  facing_item[curtain_143,drawing_140]=True
  inside[wall_26,dining_room_1]=True
  facing_item[shower_167,drawing_186]=True
  on[pot_98,oven_82]=True
  inside[wall_246,bedroom_189]=True
  inside[pillow_287,home_office_248]=True
  close_item[couch_71,powersocket_197]=True
  close_item[couch_71,floor_5]=True
  close_item[couch_71,photoframe_133]=True
  close_item[couch_71,floor_6]=True
  close_item[couch_71,orchid_136]=True
  close_item[couch_71,nightstand_72]=True
  close_item[couch_71,drawing_138]=True
  close_item[couch_71,drawing_139]=True
  close_item[couch_71,drawing_140]=True
  close_item[couch_71,drawing_141]=True
  close_item[couch_71,drawing_142]=True
  close_item[couch_71,nightstand_73]=True
  close_item[couch_71,ceiling_16]=True
  close_item[couch_71,dog_2000]=True
  close_item[couch_71,clothes_hat_2001]=True
  close_item[couch_71,clothes_hat_2028]=True
  close_item[couch_71,clothes_scarf_2004]=True
  close_item[couch_71,wall_22]=True
  close_item[couch_71,wall_23]=True
  close_item[microwave_86,cupboard_65]=True
  close_item[microwave_86,kitchen_counter_66]=True
  close_item[microwave_86,sink_67]=True
  close_item[microwave_86,faucet_68]=True
  close_item[microwave_86,floor_9]=True
  close_item[microwave_86,ceiling_13]=True
  close_item[microwave_86,food_butter_2035]=True
  close_item[microwave_86,phone_148]=True
  close_item[microwave_86,wall_21]=True
  close_item[microwave_86,wall_24]=True
  close_item[toaster_76,pot_97]=True
  close_item[toaster_76,kitchen_counter_66]=True
  close_item[toaster_76,sink_67]=True
  close_item[toaster_76,faucet_68]=True
  close_item[toaster_76,pot_98]=True
  close_item[toaster_76,walllamp_36]=True
  close_item[toaster_76,cupboard_65]=True
  close_item[toaster_76,floor_9]=True
  close_item[toaster_76,floor_11]=True
  close_item[toaster_76,ceiling_12]=True
  close_item[toaster_76,ceiling_13]=True
  close_item[toaster_76,stovefan_79]=True
  close_item[toaster_76,oven_82]=True
  close_item[toaster_76,tray_83]=True
  close_item[toaster_76,wall_21]=True
  close_item[toaster_76,wall_24]=True
  close_item[toaster_76,wall_26]=True
  close_item[toaster_76,knifeblock_92]=True
  close_item[shower_169,floor_161]=True
  close_item[shower_169,ceilinglamp_164]=True
  close_item[shower_169,photoframe_133]=True
  close_item[shower_169,toilet_166]=True
  close_item[shower_169,shower_167]=True
  close_item[shower_169,floor_6]=True
  close_item[shower_169,nightstand_73]=True
  close_item[shower_169,curtain_170]=True
  close_item[shower_169,freezer_80]=True
  close_item[shower_169,ceiling_17]=True
  close_item[shower_169,wall_22]=True
  close_item[shower_169,wall_153]=True
  close_item[shower_169,ceiling_156]=True
  inside[bed_194,bedroom_189]=True
  close_item[bookshelf_190,doorjamb_228]=True
  close_item[bookshelf_190,powersocket_197]=True
  close_item[bookshelf_190,mat_230]=True
  close_item[bookshelf_190,door_229]=True
  close_item[bookshelf_190,floor_234]=True
  close_item[bookshelf_190,floor_235]=True
  close_item[bookshelf_190,photoframe_204]=True
  close_item[bookshelf_190,floor_236]=True
  close_item[bookshelf_190,ceiling_239]=True
  close_item[bookshelf_190,ceiling_240]=True
  close_item[bookshelf_190,wall_243]=True
  close_item[bookshelf_190,wall_245]=True
  close_item[bookshelf_190,form_2015]=True
  close_item[bookshelf_190,chair_191]=True
  facing_item[ceiling_157,drawing_186]=True
  inside[ceilinglamp_35,dining_room_1]=True
  inside[floor_158,bathroom_149]=True
  facing_item[orchid_282,computer_273]=True
  facing_item[orchid_282,drawing_283]=True
  facing_item[orchid_282,television_278]=True
  close_item[ceiling_333,wall_321]=True
  close_item[ceiling_333,hanger_259]=True
  close_item[ceiling_333,hanger_260]=True
  close_item[ceiling_333,wall_324]=True
  close_item[ceiling_333,wall_325]=True
  close_item[ceiling_333,hanger_261]=True
  close_item[ceiling_333,ceiling_330]=True
  close_item[ceiling_333,ceiling_332]=True
  close_item[ceiling_333,ceiling_334]=True
  close_item[ceiling_333,television_278]=True
  close_item[ceiling_333,window_348]=True
  close_item[ceiling_333,walllamp_316]=True
  close_item[ceiling_333,walllamp_315]=True
  close_item[ceiling_333,curtain_284]=True
  close_item[ceiling_333,curtain_285]=True
  close_item[ceiling_333,curtain_286]=True
  inside[nightstand_255,home_office_248]=True
  on[tablelamp_317,nightstand_255]=True
  close_item[floor_338,desk_192]=True
  close_item[floor_338,wall_322]=True
  close_item[floor_338,filing_cabinet_195]=True
  close_item[floor_338,door_347]=True
  close_item[floor_338,floor_236]=True
  close_item[floor_338,floor_337]=True
  close_item[floor_338,cpuscreen_274]=True
  close_item[floor_338,keyboard_275]=True
  close_item[floor_338,floor_339]=True
  close_item[floor_338,computer_273]=True
  close_item[floor_338,wall_245]=True
  close_item[floor_338,walllamp_311]=True
  close_item[floor_338,light_280]=True
  close_item[floor_338,mat_281]=True
  close_item[floor_338,bookshelf_250]=True
  close_item[floor_338,desk_251]=True
  close_item[floor_338,chair_254]=True
  on[clothes_dress_2007,couch_257]=True
  on[knife_2064,mat_135]=True
  inside[ceiling_239,bedroom_189]=True
  close_item[knife_2024,cupboard_65]=True
  inside[shower_167,bathroom_149]=True
  inside[cup_1001,bedroom_189]=True
  inside[light_187,bathroom_149]=True
  on[sheets_2032,bed_194]=True
  inside[wall_151,bathroom_149]=True
  facing_item[ceiling_16,drawing_139]=True
  facing_item[ceiling_16,drawing_140]=True
  facing_item[ceiling_16,drawing_141]=True
  facing_item[ceiling_16,drawing_142]=True
  close_item[ceilinglamp_233,ceiling_239]=True
  close_item[ceilinglamp_233,ceiling_240]=True
  close_item[ceilinglamp_233,ceiling_241]=True
  close_item[ceilinglamp_233,ceiling_242]=True
  close_item[ceilinglamp_233,wall_243]=True
  close_item[ceilinglamp_233,wall_244]=True
  close_item[ceilinglamp_233,wall_245]=True
  close_item[ceilinglamp_233,wall_246]=True
  inside[floor_2,dining_room_1]=True
  inside[coffee_filter_2050,dining_room_1]=True
  on[table_63,floor_4]=True
  facing_item[floor_341,drawing_283]=True
  on[shower_169,floor_161]=True
  facing_item[closetdrawer_268,computer_273]=True
  inside[curtain_170,shower_169]=True
  inside[curtain_170,bathroom_149]=True
  on[photoframe_133,nightstand_73]=True
  facing_item[ceiling_15,drawing_139]=True
  facing_item[ceiling_15,drawing_140]=True
  facing_item[ceiling_15,drawing_141]=True
  facing_item[ceiling_15,drawing_142]=True
  inside[ceiling_154,bathroom_149]=True
  close_item[door_229,nightstand_193]=True
  close_item[door_229,doorjamb_228]=True
  close_item[door_229,powersocket_197]=True
  close_item[door_229,mat_230]=True
  close_item[door_229,floor_5]=True
  close_item[door_229,floor_8]=True
  close_item[door_229,orchid_136]=True
  close_item[door_229,floor_234]=True
  close_item[door_229,floor_235]=True
  close_item[door_229,nightstand_72]=True
  close_item[door_229,wallshelf_75]=True
  close_item[door_229,wallshelf_74]=True
  close_item[door_229,floor_238]=True
  close_item[door_229,wall_243]=True
  close_item[door_229,wall_244]=True
  close_item[door_229,wall_23]=True
  close_item[door_229,bookshelf_190]=True
  close_item[door_229,wall_30]=True
  inside[plate_1004,dishwasher_1002]=True
  inside[plate_1004,bedroom_189]=True
  close_item[floor_235,nightstand_193]=True
  close_item[floor_235,bed_194]=True
  close_item[floor_235,doorjamb_228]=True
  close_item[floor_235,door_229]=True
  close_item[floor_235,powersocket_197]=True
  close_item[floor_235,mat_230]=True
  close_item[floor_235,pillow_231]=True
  close_item[floor_235,nightstand_72]=True
  close_item[floor_235,floor_234]=True
  close_item[floor_235,orchid_136]=True
  close_item[floor_235,photoframe_204]=True
  close_item[floor_235,floor_236]=True
  close_item[floor_235,floor_238]=True
  close_item[floor_235,floor_8]=True
  close_item[floor_235,wall_243]=True
  close_item[floor_235,wall_244]=True
  close_item[floor_235,wall_245]=True
  close_item[floor_235,wall_30]=True
  close_item[floor_235,bookshelf_190]=True
  close_item[floor_235,chair_191]=True
  close_item[ceiling_240,wall_322]=True
  close_item[ceiling_240,ceiling_328]=True
  close_item[ceiling_240,ceilinglamp_233]=True
  close_item[ceiling_240,photoframe_204]=True
  close_item[ceiling_240,ceiling_239]=True
  close_item[ceiling_240,ceiling_241]=True
  close_item[ceiling_240,wall_243]=True
  close_item[ceiling_240,wall_245]=True
  close_item[ceiling_240,wall_246]=True
  close_item[ceiling_240,bookshelf_250]=True
  close_item[ceiling_240,bookshelf_190]=True
  close_item[floor_4,floor_2]=True
  close_item[floor_4,floor_3]=True
  close_item[floor_4,floor_5]=True
  close_item[floor_4,floor_7]=True
  close_item[floor_4,mat_135]=True
  close_item[floor_4,floor_11]=True
  close_item[floor_4,chair_59]=True
  close_item[floor_4,chair_60]=True
  close_item[floor_4,chair_61]=True
  close_item[floor_4,chair_62]=True
  close_item[floor_4,table_63]=True
  close_item[ceiling_19,cupboard_64]=True
  close_item[ceiling_19,ceilinglamp_35]=True
  close_item[ceiling_19,ceiling_12]=True
  close_item[ceiling_19,stovefan_79]=True
  close_item[ceiling_19,curtain_145]=True
  close_item[ceiling_19,ceiling_18]=True
  close_item[ceiling_19,coffe_maker_84]=True
  close_item[ceiling_19,wall_25]=True
  close_item[ceiling_19,wall_29]=True
  on[food_food_2031,kitchen_counter_69]=True
  close_item[clothes_socks_2052,filing_cabinet_195]=True
  close_item[wall_24,cupboard_65]=True
  close_item[wall_24,kitchen_counter_66]=True
  close_item[wall_24,sink_67]=True
  close_item[wall_24,faucet_68]=True
  close_item[wall_24,walllamp_36]=True
  close_item[wall_24,pot_98]=True
  close_item[wall_24,pot_97]=True
  close_item[wall_24,floor_9]=True
  close_item[wall_24,toaster_76]=True
  close_item[wall_24,ceiling_13]=True
  close_item[wall_24,ceiling_12]=True
  close_item[wall_24,stovefan_79]=True
  close_item[wall_24,oven_82]=True
  close_item[wall_24,tray_83]=True
  close_item[wall_24,wall_21]=True
  close_item[wall_24,microwave_86]=True
  close_item[wall_24,wall_26]=True
  close_item[wall_24,knifeblock_92]=True
  close_item[wooden_spoon_2067,kitchen_counter_70]=True
  close_item[detergent_2006,bathroom_cabinet_168]=True
  facing_item[wallshelf_75,drawing_138]=True
  facing_item[wallshelf_75,drawing_139]=True
  facing_item[wallshelf_75,drawing_140]=True
  facing_item[wallshelf_75,drawing_141]=True
  close_item[cd_2011,filing_cabinet_195]=True
  inside[wall_322,home_office_248]=True
  close_item[food_food_2031,kitchen_counter_69]=True
  close_item[pasta_2036,table_63]=True
  inside[walllamp_163,bathroom_149]=True
  close_item[hanger_262,dresser_258]=True
  close_item[hanger_262,hanger_259]=True
  close_item[hanger_262,hanger_260]=True
  close_item[hanger_262,hanger_261]=True
  close_item[hanger_262,wall_325]=True
  close_item[hanger_262,hanger_263]=True
  close_item[hanger_262,hanger_264]=True
  close_item[hanger_262,hanger_265]=True
  close_item[hanger_262,closetdrawer_266]=True
  close_item[hanger_262,closetdrawer_267]=True
  close_item[hanger_262,closetdrawer_268]=True
  close_item[hanger_262,closetdrawer_269]=True
  close_item[hanger_262,ceiling_334]=True
  close_item[hanger_262,closetdrawer_270]=True
  close_item[hanger_262,doorjamb_346]=True
  close_item[hanger_262,walllamp_315]=True
  close_item[closetdrawer_266,dresser_258]=True
  close_item[closetdrawer_266,hanger_259]=True
  close_item[closetdrawer_266,hanger_260]=True
  close_item[closetdrawer_266,wall_325]=True
  close_item[closetdrawer_266,hanger_262]=True
  close_item[closetdrawer_266,hanger_263]=True
  close_item[closetdrawer_266,hanger_261]=True
  close_item[closetdrawer_266,hanger_265]=True
  close_item[closetdrawer_266,hanger_264]=True
  close_item[closetdrawer_266,closetdrawer_267]=True
  close_item[closetdrawer_266,closetdrawer_268]=True
  close_item[closetdrawer_266,closetdrawer_269]=True
  close_item[closetdrawer_266,closetdrawer_270]=True
  close_item[closetdrawer_266,closetdrawer_271]=True
  close_item[closetdrawer_266,closetdrawer_272]=True
  close_item[closetdrawer_266,floor_344]=True
  close_item[closetdrawer_266,doorjamb_346]=True
  close_item[closetdrawer_266,walllamp_315]=True
  facing_item[ceiling_327,computer_273]=True
  facing_item[ceiling_327,drawing_283]=True
  facing_item[ceiling_154,drawing_186]=True
  close_item[mat_281,wall_320]=True
  close_item[mat_281,wall_322]=True
  close_item[mat_281,filing_cabinet_195]=True
  close_item[mat_281,light_196]=True
  close_item[mat_281,wall_323]=True
  close_item[mat_281,floor_237]=True
  close_item[mat_281,basket_for_clothes_2062]=True
  close_item[mat_281,floor_335]=True
  close_item[mat_281,floor_336]=True
  close_item[mat_281,floor_337]=True
  close_item[mat_281,floor_338]=True
  close_item[mat_281,floor_340]=True
  close_item[mat_281,wall_246]=True
  close_item[mat_281,powersocket_279]=True
  close_item[mat_281,light_280]=True
  close_item[mat_281,doorjamb_345]=True
  close_item[mat_281,bookshelf_250]=True
  close_item[mat_281,door_347]=True
  close_item[mat_281,bookshelf_253]=True
  close_item[mat_281,chair_254]=True
  close_item[pillow_287,pillow_288]=True
  close_item[pillow_287,couch_256]=True
  close_item[pillow_287,wall_324]=True
  close_item[pillow_287,floor_340]=True
  close_item[pillow_287,floor_341]=True
  close_item[pillow_287,floor_342]=True
  close_item[pillow_287,floor_343]=True
  inside[sink_173,bathroom_counter_171]=True
  inside[sink_173,bathroom_149]=True
  inside[microwave_86,dining_room_1]=True
  inside[powersocket_147,dining_room_1]=True
  on[ceiling_241,wall_246]=True
  inside[tray_2021,home_office_248]=True
  on[ceiling_334,wall_325]=True
  on[soap_2020,kitchen_counter_70]=True
  inside[ceiling_331,home_office_248]=True
  on[food_food_2008,table_249]=True
  on[nightstand_193,floor_234]=True
  on[nightstand_193,floor_235]=True
  on[orchid_282,table_249]=True
  facing_item[couch_256,television_278]=True
  close_item[table_63,ceilinglamp_34]=True
  close_item[table_63,ceilinglamp_35]=True
  close_item[table_63,floor_4]=True
  close_item[table_63,floor_5]=True
  close_item[table_63,floor_7]=True
  close_item[table_63,cutting_board_2025]=True
  close_item[table_63,floor_11]=True
  close_item[table_63,pasta_2036]=True
  close_item[table_63,chair_59]=True
  close_item[table_63,chair_60]=True
  close_item[table_63,chair_61]=True
  close_item[table_63,chair_62]=True
  inside[walllamp_315,home_office_248]=True
  close_item[plate_1005,food_food_2033]=True
  close_item[faucet_68,cupboard_65]=True
  close_item[faucet_68,kitchen_counter_66]=True
  close_item[faucet_68,sink_67]=True
  close_item[faucet_68,floor_9]=True
  close_item[faucet_68,floor_11]=True
  close_item[faucet_68,toaster_76]=True
  close_item[faucet_68,ceiling_13]=True
  close_item[faucet_68,wall_21]=True
  close_item[faucet_68,microwave_86]=True
  close_item[faucet_68,wall_24]=True
  close_item[faucet_68,wall_26]=True
  close_item[faucet_68,knifeblock_92]=True
  close_item[tray_83,cupboard_64]=True
  close_item[tray_83,pot_97]=True
  close_item[tray_83,pot_98]=True
  close_item[tray_83,kitchen_counter_66]=True
  close_item[tray_83,walllamp_36]=True
  close_item[tray_83,kitchen_counter_69]=True
  close_item[tray_83,cupboard_65]=True
  close_item[tray_83,floor_9]=True
  close_item[tray_83,floor_11]=True
  close_item[tray_83,toaster_76]=True
  close_item[tray_83,stovefan_79]=True
  close_item[tray_83,oven_82]=True
  close_item[tray_83,wall_21]=True
  close_item[tray_83,wall_24]=True
  close_item[tray_83,wall_25]=True
  close_item[tray_83,wall_26]=True
  close_item[tray_83,knifeblock_92]=True
  close_item[tray_83,wall_29]=True
  on[ceiling_157,wall_152]=True
  on[clothes_hat_2001,couch_71]=True
  inside[soap_2030,dining_room_1]=True
  inside[powersocket_279,home_office_248]=True
  close_item[pillow_288,couch_256]=True
  close_item[pillow_288,nightstand_255]=True
  close_item[pillow_288,wall_324]=True
  close_item[pillow_288,wall_323]=True
  close_item[pillow_288,floor_340]=True
  close_item[pillow_288,floor_341]=True
  close_item[pillow_288,floor_342]=True
  close_item[pillow_288,floor_343]=True
  close_item[pillow_288,table_249]=True
  close_item[pillow_288,tablelamp_317]=True
  close_item[pillow_288,pillow_287]=True
  facing_item[floor_3,drawing_138]=True
  facing_item[floor_3,drawing_139]=True
  facing_item[floor_3,drawing_140]=True
  facing_item[floor_3,drawing_141]=True
  facing_item[floor_3,drawing_142]=True
  inside[knife_2024,cupboard_65]=True
  inside[knife_2024,dining_room_1]=True
  on[toaster_76,kitchen_counter_66]=True
  close_item[wall_325,dresser_258]=True
  close_item[wall_325,hanger_259]=True
  close_item[wall_325,hanger_260]=True
  close_item[wall_325,hanger_261]=True
  close_item[wall_325,hanger_262]=True
  close_item[wall_325,hanger_263]=True
  close_item[wall_325,hanger_264]=True
  close_item[wall_325,hanger_265]=True
  close_item[wall_325,closetdrawer_266]=True
  close_item[wall_325,closetdrawer_267]=True
  close_item[wall_325,closetdrawer_268]=True
  close_item[wall_325,closetdrawer_269]=True
  close_item[wall_325,closetdrawer_270]=True
  close_item[wall_325,closetdrawer_271]=True
  close_item[wall_325,closetdrawer_272]=True
  close_item[wall_325,computer_273]=True
  close_item[wall_325,mousepad_276]=True
  close_item[wall_325,mouse_277]=True
  close_item[wall_325,television_278]=True
  close_item[wall_325,curtain_284]=True
  close_item[wall_325,curtain_285]=True
  close_item[wall_325,walllamp_312]=True
  close_item[wall_325,walllamp_315]=True
  close_item[wall_325,wall_319]=True
  close_item[wall_325,wall_321]=True
  close_item[wall_325,ceiling_329]=True
  close_item[wall_325,ceiling_333]=True
  close_item[wall_325,ceiling_334]=True
  close_item[wall_325,floor_339]=True
  close_item[wall_325,floor_343]=True
  close_item[wall_325,floor_344]=True
  close_item[wall_325,doorjamb_346]=True
  close_item[wall_325,window_348]=True
  close_item[wall_325,tvstand_252]=True
  on[cupboard_64,wall_29]=True
  close_item[doorjamb_345,wall_320]=True
  close_item[doorjamb_345,wall_322]=True
  close_item[doorjamb_345,filing_cabinet_195]=True
  close_item[doorjamb_345,light_196]=True
  close_item[doorjamb_345,wall_323]=True
  close_item[doorjamb_345,ceiling_327]=True
  close_item[doorjamb_345,floor_237]=True
  close_item[doorjamb_345,floor_337]=True
  close_item[doorjamb_345,ceiling_241]=True
  close_item[doorjamb_345,wall_245]=True
  close_item[doorjamb_345,wall_246]=True
  close_item[doorjamb_345,powersocket_279]=True
  close_item[doorjamb_345,light_280]=True
  close_item[doorjamb_345,mat_281]=True
  close_item[doorjamb_345,bookshelf_250]=True
  close_item[doorjamb_345,door_347]=True
  close_item[doorjamb_345,bookshelf_253]=True
  between[door_347,home_office_248]=True
  between[door_347,bedroom_189]=True
  facing_item[table_249,computer_273]=True
  facing_item[table_249,drawing_283]=True
  facing_item[table_249,television_278]=True
  inside[ceiling_334,home_office_248]=True
  facing_item[powersocket_279,drawing_283]=True
  inside[pot_98,dining_room_1]=True
  facing_item[ceiling_17,drawing_139]=True
  facing_item[ceiling_17,drawing_140]=True
  facing_item[ceiling_17,drawing_141]=True
  facing_item[ceiling_17,drawing_142]=True
  close_item[dishwasher_81,cupboard_64]=True
  close_item[dishwasher_81,pot_97]=True
  close_item[dishwasher_81,pot_98]=True
  close_item[dishwasher_81,kitchen_counter_69]=True
  close_item[dishwasher_81,kitchen_counter_70]=True
  close_item[dishwasher_81,floor_10]=True
  close_item[dishwasher_81,floor_11]=True
  close_item[dishwasher_81,coffe_maker_84]=True
  close_item[dishwasher_81,wall_25]=True
  close_item[dishwasher_81,wall_26]=True
  close_item[dishwasher_81,wall_29]=True
  close_item[bathroom_cabinet_168,walllamp_163]=True
  close_item[bathroom_cabinet_168,walllamp_165]=True
  close_item[bathroom_cabinet_168,bathroom_counter_171]=True
  close_item[bathroom_cabinet_168,faucet_172]=True
  close_item[bathroom_cabinet_168,sink_173]=True
  close_item[bathroom_cabinet_168,detergent_2006]=True
  close_item[bathroom_cabinet_168,wall_151]=True
  close_item[bathroom_cabinet_168,wall_152]=True
  close_item[bathroom_cabinet_168,ceiling_154]=True
  close_item[bathroom_cabinet_168,ceiling_157]=True
  inside[orchid_282,home_office_248]=True
  inside[food_food_2033,bedroom_189]=True
  facing_item[walllamp_315,computer_273]=True
  facing_item[floor_158,drawing_186]=True
  inside[chair_62,dining_room_1]=True
  close_item[knife_2064,mat_135]=True
  on[keyboard_2057,desk_251]=True
  inside[knife_2017,bedroom_189]=True
  close_item[ceiling_332,pillow_289]=True
  close_item[ceiling_332,couch_257]=True
  close_item[ceiling_332,wall_324]=True
  close_item[ceiling_332,ceiling_331]=True
  close_item[ceiling_332,ceiling_333]=True
  close_item[ceiling_332,walllamp_316]=True
  close_item[ceiling_332,curtain_286]=True
  close_item[door_347,wall_320]=True
  close_item[door_347,wall_322]=True
  close_item[door_347,filing_cabinet_195]=True
  close_item[door_347,light_196]=True
  close_item[door_347,wall_323]=True
  close_item[door_347,mat_281]=True
  close_item[door_347,floor_236]=True
  close_item[door_347,floor_237]=True
  close_item[door_347,floor_335]=True
  close_item[door_347,floor_336]=True
  close_item[door_347,floor_337]=True
  close_item[door_347,floor_338]=True
  close_item[door_347,wall_245]=True
  close_item[door_347,wall_246]=True
  close_item[door_347,powersocket_279]=True
  close_item[door_347,light_280]=True
  close_item[door_347,doorjamb_345]=True
  close_item[door_347,bookshelf_250]=True
  close_item[door_347,bookshelf_253]=True
  inside[floor_343,home_office_248]=True
  on[door_229,floor_234]=True
  on[door_229,floor_235]=True
  close_item[wall_29,floor_7]=True
  close_item[wall_29,floor_10]=True
  close_item[wall_29,floor_11]=True
  close_item[wall_29,ceiling_12]=True
  close_item[wall_29,curtain_145]=True
  close_item[wall_29,ceiling_18]=True
  close_item[wall_29,ceiling_19]=True
  close_item[wall_29,wall_25]=True
  close_item[wall_29,wall_26]=True
  close_item[wall_29,wall_27]=True
  close_item[wall_29,window_33]=True
  close_item[wall_29,ceilinglamp_35]=True
  close_item[wall_29,walllamp_36]=True
  close_item[wall_29,chair_62]=True
  close_item[wall_29,cupboard_64]=True
  close_item[wall_29,kitchen_counter_69]=True
  close_item[wall_29,kitchen_counter_70]=True
  close_item[wall_29,stovefan_79]=True
  close_item[wall_29,dishwasher_81]=True
  close_item[wall_29,oven_82]=True
  close_item[wall_29,tray_83]=True
  close_item[wall_29,coffe_maker_84]=True
  close_item[wall_29,pot_97]=True
  close_item[wall_29,pot_98]=True
  close_item[ceilinglamp_34,ceiling_12]=True
  close_item[ceilinglamp_34,ceiling_13]=True
  close_item[ceilinglamp_34,ceiling_14]=True
  close_item[ceilinglamp_34,ceiling_15]=True
  close_item[ceilinglamp_34,ceiling_16]=True
  close_item[ceilinglamp_34,ceiling_17]=True
  close_item[ceilinglamp_34,wall_21]=True
  close_item[ceilinglamp_34,wall_22]=True
  close_item[ceilinglamp_34,chair_59]=True
  close_item[ceilinglamp_34,chair_61]=True
  close_item[ceilinglamp_34,table_63]=True
  facing_item[nightstand_72,drawing_140]=True
  inside[floor_337,home_office_248]=True
  inside[bookshelf_250,home_office_248]=True
  on[cutting_board_2025,table_63]=True
  inside[cupboard_65,dining_room_1]=True
  inside[keyboard_275,home_office_248]=True
  facing_item[wall_324,drawing_283]=True
  facing_item[wall_324,television_278]=True
  inside[dog_2000,dining_room_1]=True
  facing_item[window_348,television_278]=True
  inside[pasta_2036,dining_room_1]=True
  inside[wall_29,dining_room_1]=True
  close_item[pillow_232,bed_194]=True
  close_item[pillow_232,wall_244]=True
  close_item[pillow_232,floor_238]=True
  close_item[pillow_232,pillow_231]=True
  inside[doorjamb_346,home_office_248]=True
  inside[ceiling_13,dining_room_1]=True
  inside[ceilinglamp_310,home_office_248]=True
  close_item[check_2003,couch_256]=True
  inside[toothbrush_holder_2061,bathroom_149]=True
  close_item[mat_135,doorjamb_32]=True
  close_item[mat_135,floor_160]=True
  close_item[mat_135,floor_2]=True
  close_item[mat_135,floor_3]=True
  close_item[mat_135,floor_4]=True
  close_item[mat_135,toilet_166]=True
  close_item[mat_135,floor_6]=True
  close_item[mat_135,shower_167]=True
  close_item[mat_135,floor_9]=True
  close_item[mat_135,freezer_80]=True
  close_item[mat_135,knife_2064]=True
  close_item[mat_135,light_146]=True
  close_item[mat_135,powersocket_147]=True
  close_item[mat_135,wall_21]=True
  close_item[mat_135,wall_150]=True
  close_item[mat_135,wall_22]=True
  close_item[mat_135,light_187]=True
  close_item[mat_135,wall_28]=True
  close_item[mat_135,door_31]=True
  on[dishwasher_81,floor_10]=True
  close_item[wall_150,floor_2]=True
  close_item[wall_150,floor_3]=True
  close_item[wall_150,mat_135]=True
  close_item[wall_150,ceiling_14]=True
  close_item[wall_150,light_146]=True
  close_item[wall_150,powersocket_147]=True
  close_item[wall_150,phone_148]=True
  close_item[wall_150,wall_151]=True
  close_item[wall_150,wall_153]=True
  close_item[wall_150,ceiling_154]=True
  close_item[wall_150,ceiling_155]=True
  close_item[wall_150,ceiling_156]=True
  close_item[wall_150,wall_28]=True
  close_item[wall_150,floor_158]=True
  close_item[wall_150,floor_159]=True
  close_item[wall_150,floor_160]=True
  close_item[wall_150,doorjamb_32]=True
  close_item[wall_150,floor_161]=True
  close_item[wall_150,door_31]=True
  close_item[wall_150,ceilinglamp_164]=True
  close_item[wall_150,toilet_166]=True
  close_item[wall_150,shower_167]=True
  close_item[wall_150,curtain_170]=True
  close_item[wall_150,mat_185]=True
  close_item[wall_150,light_187]=True
  close_item[wall_150,freezer_80]=True
  between[door_31,dining_room_1]=True
  between[door_31,bathroom_149]=True
  close_item[drawing_140,couch_71]=True
  close_item[drawing_140,drawing_138]=True
  close_item[drawing_140,drawing_139]=True
  close_item[drawing_140,drawing_141]=True
  close_item[drawing_140,drawing_142]=True
  close_item[drawing_140,ceiling_239]=True
  close_item[drawing_140,ceiling_16]=True
  close_item[drawing_140,ceiling_17]=True
  close_item[drawing_140,wall_243]=True
  close_item[drawing_140,ceiling_20]=True
  close_item[drawing_140,wall_22]=True
  close_item[drawing_140,wall_23]=True
  close_item[drawing_140,wall_30]=True
  close_item[ceiling_155,doorjamb_32]=True
  close_item[ceiling_155,ceilinglamp_164]=True
  close_item[ceiling_155,shower_167]=True
  close_item[ceiling_155,ceiling_14]=True
  close_item[ceiling_155,ceiling_156]=True
  close_item[ceiling_155,light_146]=True
  close_item[ceiling_155,phone_148]=True
  close_item[ceiling_155,wall_150]=True
  close_item[ceiling_155,wall_151]=True
  close_item[ceiling_155,wall_153]=True
  close_item[ceiling_155,ceiling_154]=True
  close_item[ceiling_155,light_187]=True
  close_item[ceiling_155,wall_28]=True
  inside[dresser_258,home_office_248]=True
  close_item[bookmark_2046,filing_cabinet_195]=True
  inside[food_food_2045,bedroom_189]=True
  inside[photoframe_294,home_office_248]=True
  inside[photoframe_294,bookshelf_253]=True
  facing_item[couch_257,television_278]=True
  inside[faucet_68,dining_room_1]=True
  inside[wall_22,dining_room_1]=True
  on[bookshelf_253,floor_336]=True
  on[bookshelf_253,floor_335]=True
  inside[ceiling_16,dining_room_1]=True
  facing_item[wall_151,drawing_186]=True
  inside[knife_2064,dining_room_1]=True
  close_item[wall_30,floor_5]=True
  close_item[wall_30,floor_7]=True
  close_item[wall_30,floor_8]=True
  close_item[wall_30,orchid_136]=True
  close_item[wall_30,drawing_138]=True
  close_item[wall_30,drawing_140]=True
  close_item[wall_30,curtain_143]=True
  close_item[wall_30,curtain_144]=True
  close_item[wall_30,ceiling_16]=True
  close_item[wall_30,ceiling_18]=True
  close_item[wall_30,ceiling_20]=True
  close_item[wall_30,wall_23]=True
  close_item[wall_30,wall_27]=True
  close_item[wall_30,window_33]=True
  close_item[wall_30,ceilinglamp_35]=True
  close_item[wall_30,chair_59]=True
  close_item[wall_30,chair_60]=True
  close_item[wall_30,nightstand_193]=True
  close_item[wall_30,powersocket_197]=True
  close_item[wall_30,nightstand_72]=True
  close_item[wall_30,wallshelf_74]=True
  close_item[wall_30,wallshelf_75]=True
  close_item[wall_30,doorjamb_228]=True
  close_item[wall_30,door_229]=True
  close_item[wall_30,pillow_231]=True
  close_item[wall_30,floor_234]=True
  close_item[wall_30,floor_235]=True
  close_item[wall_30,ceiling_239]=True
  close_item[wall_30,wall_243]=True
  facing_item[walllamp_163,drawing_186]=True
  close_item[ceilinglamp_35,ceiling_12]=True
  close_item[ceilinglamp_35,ceiling_15]=True
  close_item[ceilinglamp_35,ceiling_16]=True
  close_item[ceilinglamp_35,ceiling_18]=True
  close_item[ceilinglamp_35,ceiling_19]=True
  close_item[ceilinglamp_35,ceiling_20]=True
  close_item[ceilinglamp_35,wall_30]=True
  close_item[ceilinglamp_35,chair_60]=True
  close_item[ceilinglamp_35,wall_29]=True
  close_item[ceilinglamp_35,chair_62]=True
  close_item[ceilinglamp_35,table_63]=True
  inside[floor_236,bedroom_189]=True
  facing_item[wall_30,drawing_139]=True
  facing_item[wall_30,drawing_140]=True
  facing_item[wall_30,drawing_141]=True
  facing_item[wall_30,drawing_142]=True
  close_item[detergent_2041,filing_cabinet_195]=True
  on[shoe_rack_2013,mat_230]=True
  close_item[nightstand_193,bed_194]=True
  close_item[nightstand_193,doorjamb_228]=True
  close_item[nightstand_193,door_229]=True
  close_item[nightstand_193,powersocket_197]=True
  close_item[nightstand_193,pillow_231]=True
  close_item[nightstand_193,mat_230]=True
  close_item[nightstand_193,floor_8]=True
  close_item[nightstand_193,floor_234]=True
  close_item[nightstand_193,floor_235]=True
  close_item[nightstand_193,floor_238]=True
  close_item[nightstand_193,wall_243]=True
  close_item[nightstand_193,wall_244]=True
  close_item[nightstand_193,wall_30]=True
  close_item[light_280,wall_320]=True
  close_item[light_280,desk_192]=True
  close_item[light_280,wall_322]=True
  close_item[light_280,filing_cabinet_195]=True
  close_item[light_280,light_196]=True
  close_item[light_280,mat_281]=True
  close_item[light_280,ceiling_327]=True
  close_item[light_280,floor_236]=True
  close_item[light_280,floor_237]=True
  close_item[light_280,floor_337]=True
  close_item[light_280,ceiling_241]=True
  close_item[light_280,floor_338]=True
  close_item[light_280,wall_245]=True
  close_item[light_280,wall_246]=True
  close_item[light_280,powersocket_279]=True
  close_item[light_280,doorjamb_345]=True
  close_item[light_280,bookshelf_250]=True
  close_item[light_280,door_347]=True
  inside[thread_2012,filing_cabinet_195]=True
  inside[thread_2012,bedroom_189]=True
  inside[hanger_261,home_office_248]=True
  inside[hanger_261,dresser_258]=True
  inside[wall_25,dining_room_1]=True
  close_item[ceiling_239,doorjamb_228]=True
  close_item[ceiling_239,ceilinglamp_233]=True
  close_item[ceiling_239,drawing_138]=True
  close_item[ceiling_239,photoframe_204]=True
  close_item[ceiling_239,drawing_140]=True
  close_item[ceiling_239,ceiling_240]=True
  close_item[ceiling_239,ceiling_242]=True
  close_item[ceiling_239,wall_243]=True
  close_item[ceiling_239,ceiling_20]=True
  close_item[ceiling_239,wall_244]=True
  close_item[ceiling_239,wall_245]=True
  close_item[ceiling_239,wall_30]=True
  close_item[ceiling_239,bookshelf_190]=True
  on[ceiling_242,wall_244]=True
  facing_item[pillow_290,television_278]=True
  inside[wall_245,bedroom_189]=True
  facing_item[wall_318,television_278]=True
  inside[floor_9,dining_room_1]=True
  inside[keyboard_2057,home_office_248]=True
  close_item[check_2002,bookshelf_253]=True
  close_item[knife_2017,kitchen_counter_1000]=True
  inside[nightstand_193,bedroom_189]=True
  inside[door_229,bedroom_189]=True
  inside[closetdrawer_270,home_office_248]=True
  inside[closetdrawer_270,dresser_258]=True
  on[kitchen_counter_69,floor_10]=True
  close_item[nightstand_73,floor_161]=True
  close_item[nightstand_73,photoframe_133]=True
  close_item[nightstand_73,floor_6]=True
  close_item[nightstand_73,couch_71]=True
  close_item[nightstand_73,floor_5]=True
  close_item[nightstand_73,shower_169]=True
  close_item[nightstand_73,drawing_142]=True
  close_item[nightstand_73,freezer_80]=True
  close_item[nightstand_73,wall_22]=True
  close_item[nightstand_73,wall_23]=True
  close_item[nightstand_73,wall_153]=True
  close_item[plate_1004,food_carrot_2018]=True
  close_item[plate_1004,food_food_2045]=True
  close_item[food_orange_2042,freezer_80]=True
  on[check_2002,bookshelf_253]=True
  facing_item[nightstand_73,drawing_141]=True
  facing_item[nightstand_73,drawing_142]=True
  close_item[floor_237,wall_320]=True
  close_item[floor_237,desk_192]=True
  close_item[floor_237,bed_194]=True
  close_item[floor_237,filing_cabinet_195]=True
  close_item[floor_237,light_196]=True
  close_item[floor_237,mat_281]=True
  close_item[floor_237,mat_230]=True
  close_item[floor_237,floor_236]=True
  close_item[floor_237,floor_238]=True
  close_item[floor_237,floor_337]=True
  close_item[floor_237,wall_244]=True
  close_item[floor_237,wall_245]=True
  close_item[floor_237,wall_246]=True
  close_item[floor_237,powersocket_279]=True
  close_item[floor_237,light_280]=True
  close_item[floor_237,doorjamb_345]=True
  close_item[floor_237,bookshelf_250]=True
  close_item[floor_237,door_347]=True
  close_item[floor_237,bookshelf_253]=True
  inside[drawing_141,dining_room_1]=True
  close_item[wall_324,couch_256]=True
  close_item[wall_324,couch_257]=True
  close_item[wall_324,orchid_282]=True
  close_item[wall_324,curtain_286]=True
  close_item[wall_324,pillow_287]=True
  close_item[wall_324,pillow_288]=True
  close_item[wall_324,pillow_289]=True
  close_item[wall_324,pillow_290]=True
  close_item[wall_324,walllamp_316]=True
  close_item[wall_324,tablelamp_317]=True
  close_item[wall_324,wall_318]=True
  close_item[wall_324,wall_321]=True
  close_item[wall_324,ceiling_331]=True
  close_item[wall_324,ceiling_332]=True
  close_item[wall_324,ceiling_333]=True
  close_item[wall_324,floor_341]=True
  close_item[wall_324,floor_342]=True
  close_item[wall_324,floor_343]=True
  close_item[wall_324,window_348]=True
  close_item[wall_324,table_249]=True
  close_item[wall_324,nightstand_255]=True
  close_item[floor_339,wall_322]=True
  close_item[floor_339,floor_344]=True
  close_item[floor_339,wall_325]=True
  close_item[floor_339,computer_273]=True
  close_item[floor_339,cpuscreen_274]=True
  close_item[floor_339,keyboard_275]=True
  close_item[floor_339,mousepad_276]=True
  close_item[floor_339,mouse_277]=True
  close_item[floor_339,floor_340]=True
  close_item[floor_339,floor_338]=True
  close_item[floor_339,walllamp_312]=True
  close_item[floor_339,television_278]=True
  close_item[floor_339,desk_251]=True
  close_item[floor_339,tvstand_252]=True
  close_item[floor_339,chair_254]=True
  close_item[floor_339,wall_319]=True
  close_item[clothes_underwear_2049,couch_257]=True
  close_item[floor_344,dresser_258]=True
  close_item[floor_344,wall_325]=True
  close_item[floor_344,closetdrawer_266]=True
  close_item[floor_344,closetdrawer_267]=True
  close_item[floor_344,closetdrawer_268]=True
  close_item[floor_344,closetdrawer_269]=True
  close_item[floor_344,closetdrawer_270]=True
  close_item[floor_344,closetdrawer_271]=True
  close_item[floor_344,closetdrawer_272]=True
  close_item[floor_344,computer_273]=True
  close_item[floor_344,floor_339]=True
  close_item[floor_344,mouse_277]=True
  close_item[floor_344,television_278]=True
  close_item[floor_344,floor_343]=True
  close_item[floor_344,doorjamb_346]=True
  close_item[floor_344,walllamp_315]=True
  close_item[floor_344,tvstand_252]=True
  close_item[wall_21,floor_2]=True
  close_item[wall_21,floor_3]=True
  close_item[wall_21,mat_135]=True
  close_item[wall_21,floor_9]=True
  close_item[wall_21,floor_11]=True
  close_item[wall_21,ceiling_12]=True
  close_item[wall_21,ceiling_13]=True
  close_item[wall_21,ceiling_14]=True
  close_item[wall_21,phone_148]=True
  close_item[wall_21,wall_24]=True
  close_item[wall_21,wall_26]=True
  close_item[wall_21,wall_28]=True
  close_item[wall_21,door_31]=True
  close_item[wall_21,doorjamb_32]=True
  close_item[wall_21,ceilinglamp_34]=True
  close_item[wall_21,walllamp_36]=True
  close_item[wall_21,light_187]=True
  close_item[wall_21,chair_61]=True
  close_item[wall_21,cupboard_65]=True
  close_item[wall_21,kitchen_counter_66]=True
  close_item[wall_21,sink_67]=True
  close_item[wall_21,faucet_68]=True
  close_item[wall_21,toaster_76]=True
  close_item[wall_21,stovefan_79]=True
  close_item[wall_21,oven_82]=True
  close_item[wall_21,tray_83]=True
  close_item[wall_21,microwave_86]=True
  close_item[wall_21,knifeblock_92]=True
  close_item[wall_21,pot_97]=True
  close_item[wall_21,pot_98]=True
  inside[floor_238,bedroom_189]=True
  close_item[wall_26,floor_11]=True
  close_item[wall_26,ceiling_12]=True
  close_item[wall_26,wall_21]=True
  close_item[wall_26,wall_24]=True
  close_item[wall_26,wall_25]=True
  close_item[wall_26,wall_29]=True
  close_item[wall_26,walllamp_36]=True
  close_item[wall_26,cupboard_64]=True
  close_item[wall_26,cupboard_65]=True
  close_item[wall_26,kitchen_counter_66]=True
  close_item[wall_26,sink_67]=True
  close_item[wall_26,faucet_68]=True
  close_item[wall_26,kitchen_counter_69]=True
  close_item[wall_26,toaster_76]=True
  close_item[wall_26,stovefan_79]=True
  close_item[wall_26,dishwasher_81]=True
  close_item[wall_26,oven_82]=True
  close_item[wall_26,tray_83]=True
  close_item[wall_26,coffe_maker_84]=True
  close_item[wall_26,knifeblock_92]=True
  close_item[wall_26,pot_97]=True
  close_item[wall_26,pot_98]=True
  inside[pillow_232,bedroom_189]=True
  inside[drawing_186,bathroom_149]=True
  on[ceiling_332,wall_324]=True
  close_item[wallshelf_74,window_33]=True
  close_item[wallshelf_74,door_229]=True
  close_item[wallshelf_74,wallshelf_75]=True
  close_item[wallshelf_74,curtain_143]=True
  close_item[wallshelf_74,curtain_144]=True
  close_item[wallshelf_74,ceiling_18]=True
  close_item[wallshelf_74,ceiling_20]=True
  close_item[wallshelf_74,wall_27]=True
  close_item[wallshelf_74,wall_30]=True
  close_item[freezer_80,floor_2]=True
  close_item[freezer_80,floor_3]=True
  close_item[freezer_80,photoframe_133]=True
  close_item[freezer_80,floor_6]=True
  close_item[freezer_80,mat_135]=True
  close_item[freezer_80,ceiling_14]=True
  close_item[freezer_80,ceiling_17]=True
  close_item[freezer_80,light_146]=True
  close_item[freezer_80,powersocket_147]=True
  close_item[freezer_80,wall_22]=True
  close_item[freezer_80,wall_150]=True
  close_item[freezer_80,wall_153]=True
  close_item[freezer_80,wall_28]=True
  close_item[freezer_80,door_31]=True
  close_item[freezer_80,doorjamb_32]=True
  close_item[freezer_80,floor_161]=True
  close_item[freezer_80,floor_160]=True
  close_item[freezer_80,toilet_166]=True
  close_item[freezer_80,shower_167]=True
  close_item[freezer_80,shower_169]=True
  close_item[freezer_80,nightstand_73]=True
  close_item[freezer_80,food_carrot_2023]=True
  close_item[freezer_80,food_orange_2042]=True
  inside[light_196,bedroom_189]=True
  inside[wall_150,bathroom_149]=True
  facing_item[nightstand_255,drawing_283]=True
  facing_item[nightstand_255,television_278]=True
  on[filing_cabinet_195,floor_237]=True
  inside[curtain_144,dining_room_1]=True
  inside[curtain_144,curtain_143]=True
  on[basket_for_clothes_2062,mat_281]=True
  facing_item[ceilinglamp_35,drawing_138]=True
  facing_item[ceilinglamp_35,drawing_139]=True
  facing_item[ceilinglamp_35,drawing_140]=True
  facing_item[ceilinglamp_35,drawing_141]=True
  facing_item[ceilinglamp_35,drawing_142]=True
  inside[ceiling_241,bedroom_189]=True
  close_item[wall_28,doorjamb_32]=True
  close_item[wall_28,floor_160]=True
  close_item[wall_28,floor_2]=True
  close_item[wall_28,floor_3]=True
  close_item[wall_28,toilet_166]=True
  close_item[wall_28,shower_167]=True
  close_item[wall_28,mat_135]=True
  close_item[wall_28,ceiling_155]=True
  close_item[wall_28,ceiling_14]=True
  close_item[wall_28,freezer_80]=True
  close_item[wall_28,light_146]=True
  close_item[wall_28,powersocket_147]=True
  close_item[wall_28,phone_148]=True
  close_item[wall_28,wall_21]=True
  close_item[wall_28,wall_150]=True
  close_item[wall_28,wall_22]=True
  close_item[wall_28,wall_153]=True
  close_item[wall_28,light_187]=True
  close_item[wall_28,door_31]=True
  close_item[drawing_142,photoframe_133]=True
  close_item[drawing_142,couch_71]=True
  close_item[drawing_142,nightstand_73]=True
  close_item[drawing_142,drawing_139]=True
  close_item[drawing_142,drawing_140]=True
  close_item[drawing_142,drawing_141]=True
  close_item[drawing_142,ceiling_16]=True
  close_item[drawing_142,ceiling_17]=True
  close_item[drawing_142,wall_22]=True
  close_item[drawing_142,wall_23]=True
  close_item[powersocket_147,doorjamb_32]=True
  close_item[powersocket_147,floor_160]=True
  close_item[powersocket_147,floor_2]=True
  close_item[powersocket_147,floor_3]=True
  close_item[powersocket_147,floor_161]=True
  close_item[powersocket_147,toilet_166]=True
  close_item[powersocket_147,mat_135]=True
  close_item[powersocket_147,shower_167]=True
  close_item[powersocket_147,floor_6]=True
  close_item[powersocket_147,freezer_80]=True
  close_item[powersocket_147,light_146]=True
  close_item[powersocket_147,wall_150]=True
  close_item[powersocket_147,wall_22]=True
  close_item[powersocket_147,wall_153]=True
  close_item[powersocket_147,wall_28]=True
  close_item[powersocket_147,door_31]=True
  facing_item[pillow_287,computer_273]=True
  facing_item[pillow_287,drawing_283]=True
  facing_item[pillow_287,television_278]=True
  on[soap_2030,kitchen_counter_70]=True
  inside[wall_153,bathroom_149]=True
  inside[cup_1003,dishwasher_1002]=True
  inside[cup_1003,bedroom_189]=True
  close_item[pillow_290,couch_257]=True
  close_item[pillow_290,pillow_289]=True
  close_item[pillow_290,wall_324]=True
  close_item[pillow_290,floor_342]=True
  close_item[pillow_290,table_249]=True
  close_item[pillow_290,walllamp_316]=True
  facing_item[floor_162,drawing_186]=True
  close_item[walllamp_311,wall_322]=True
  close_item[walllamp_311,ceiling_328]=True
  close_item[walllamp_311,ceiling_329]=True
  close_item[walllamp_311,cpuscreen_274]=True
  close_item[walllamp_311,keyboard_275]=True
  close_item[walllamp_311,floor_338]=True
  close_item[walllamp_311,desk_251]=True
  close_item[walllamp_311,wall_319]=True
  on[orchid_136,nightstand_72]=True
  on[microwave_86,kitchen_counter_66]=True
  close_item[curtain_145,window_33]=True
  close_item[curtain_145,floor_7]=True
  close_item[curtain_145,curtain_143]=True
  close_item[curtain_145,curtain_144]=True
  close_item[curtain_145,ceiling_18]=True
  close_item[curtain_145,ceiling_19]=True
  close_item[curtain_145,wall_27]=True
  close_item[curtain_145,wall_29]=True
  inside[faucet_172,bathroom_149]=True
  on[pillow_231,bed_194]=True
  close_item[knifeblock_92,cupboard_65]=True
  close_item[knifeblock_92,pot_98]=True
  close_item[knifeblock_92,sink_67]=True
  close_item[knifeblock_92,walllamp_36]=True
  close_item[knifeblock_92,faucet_68]=True
  close_item[knifeblock_92,kitchen_counter_66]=True
  close_item[knifeblock_92,pot_97]=True
  close_item[knifeblock_92,toaster_76]=True
  close_item[knifeblock_92,ceiling_12]=True
  close_item[knifeblock_92,ceiling_13]=True
  close_item[knifeblock_92,stovefan_79]=True
  close_item[knifeblock_92,oven_82]=True
  close_item[knifeblock_92,tray_83]=True
  close_item[knifeblock_92,wall_21]=True
  close_item[knifeblock_92,wall_24]=True
  close_item[knifeblock_92,wall_26]=True
  close_item[curtain_170,floor_161]=True
  close_item[curtain_170,ceilinglamp_164]=True
  close_item[curtain_170,toilet_166]=True
  close_item[curtain_170,shower_167]=True
  close_item[curtain_170,shower_169]=True
  close_item[curtain_170,wall_150]=True
  close_item[curtain_170,wall_152]=True
  close_item[curtain_170,wall_153]=True
  close_item[curtain_170,ceiling_156]=True
  close_item[mat_185,floor_160]=True
  close_item[mat_185,floor_161]=True
  close_item[mat_185,floor_162]=True
  close_item[mat_185,bathroom_counter_171]=True
  close_item[mat_185,faucet_172]=True
  close_item[mat_185,sink_173]=True
  close_item[mat_185,wall_150]=True
  close_item[mat_185,wall_151]=True
  close_item[mat_185,wall_152]=True
  close_item[mat_185,wall_153]=True
  close_item[mat_185,floor_158]=True
  close_item[mat_185,floor_159]=True
  inside[sponge_2040,bathroom_149]=True
  inside[ceiling_156,bathroom_149]=True
  close_item[chair_254,couch_256]=True
  close_item[chair_254,wall_322]=True
  close_item[chair_254,computer_273]=True
  close_item[chair_254,cpuscreen_274]=True
  close_item[chair_254,keyboard_275]=True
  close_item[chair_254,floor_339]=True
  close_item[chair_254,mousepad_276]=True
  close_item[chair_254,floor_340]=True
  close_item[chair_254,mouse_277]=True
  close_item[chair_254,floor_338]=True
  close_item[chair_254,mat_281]=True
  close_item[chair_254,floor_337]=True
  close_item[chair_254,desk_251]=True
  inside[clothes_scarf_2004,dining_room_1]=True
  inside[walllamp_314,home_office_248]=True
  close_item[needle_2009,filing_cabinet_195]=True
  close_item[dog_2000,couch_71]=True
  inside[wall_324,home_office_248]=True
  close_item[drawing_141,couch_71]=True
  close_item[drawing_141,drawing_138]=True
  close_item[drawing_141,drawing_139]=True
  close_item[drawing_141,drawing_140]=True
  close_item[drawing_141,drawing_142]=True
  close_item[drawing_141,ceiling_16]=True
  close_item[drawing_141,ceiling_17]=True
  close_item[drawing_141,wall_22]=True
  close_item[drawing_141,wall_23]=True
  close_item[light_146,floor_2]=True
  close_item[light_146,floor_3]=True
  close_item[light_146,floor_6]=True
  close_item[light_146,mat_135]=True
  close_item[light_146,ceiling_14]=True
  close_item[light_146,ceiling_17]=True
  close_item[light_146,powersocket_147]=True
  close_item[light_146,wall_150]=True
  close_item[light_146,wall_22]=True
  close_item[light_146,wall_153]=True
  close_item[light_146,ceiling_155]=True
  close_item[light_146,ceiling_156]=True
  close_item[light_146,wall_28]=True
  close_item[light_146,door_31]=True
  close_item[light_146,doorjamb_32]=True
  close_item[light_146,floor_160]=True
  close_item[light_146,floor_161]=True
  close_item[light_146,toilet_166]=True
  close_item[light_146,shower_167]=True
  close_item[light_146,light_187]=True
  close_item[light_146,freezer_80]=True
  close_item[sponge_2040,bathroom_counter_171]=True
  inside[walllamp_165,bathroom_149]=True
  inside[pencil_2039,home_office_248]=True
  inside[closetdrawer_272,home_office_248]=True
  inside[closetdrawer_272,dresser_258]=True
  close_item[desk_192,wall_322]=True
  close_item[desk_192,filing_cabinet_195]=True
  close_item[desk_192,bookmark_2053]=True
  close_item[desk_192,mat_230]=True
  close_item[desk_192,floor_236]=True
  close_item[desk_192,photoframe_204]=True
  close_item[desk_192,floor_237]=True
  close_item[desk_192,floor_338]=True
  close_item[desk_192,wall_245]=True
  close_item[desk_192,wall_246]=True
  close_item[desk_192,light_280]=True
  close_item[desk_192,bookshelf_250]=True
  close_item[desk_192,chair_191]=True
  facing_item[toilet_166,drawing_186]=True
  inside[nightstand_72,dining_room_1]=True
  on[faucet_172,bathroom_counter_171]=True
  facing_item[ceiling_20,drawing_139]=True
  facing_item[ceiling_20,drawing_140]=True
  facing_item[ceiling_20,drawing_141]=True
  facing_item[ceiling_20,drawing_142]=True
  inside[food_carrot_2023,freezer_80]=True
  inside[food_carrot_2023,dining_room_1]=True
  close_item[table_249,pillow_288]=True
  close_item[table_249,couch_257]=True
  close_item[table_249,pillow_290]=True
  close_item[table_249,wall_321]=True
  close_item[table_249,wall_324]=True
  close_item[table_249,pencil_2039]=True
  close_item[table_249,floor_340]=True
  close_item[table_249,floor_341]=True
  close_item[table_249,television_278]=True
  close_item[table_249,floor_342]=True
  close_item[table_249,walllamp_316]=True
  close_item[table_249,food_food_2008]=True
  close_item[table_249,orchid_282]=True
  close_item[table_249,dvd_player_2047]=True
  close_item[table_249,tvstand_252]=True
  close_item[table_249,floor_343]=True
  close_item[table_249,curtain_286]=True
  inside[walllamp_36,dining_room_1]=True
  inside[ceiling_333,home_office_248]=True
  facing_item[freezer_80,drawing_138]=True
  facing_item[freezer_80,drawing_139]=True
  facing_item[freezer_80,drawing_140]=True
  facing_item[freezer_80,drawing_141]=True
  facing_item[freezer_80,drawing_142]=True
  inside[mat_281,home_office_248]=True
  close_item[ceiling_157,ceilinglamp_164]=True
  close_item[ceiling_157,walllamp_165]=True
  close_item[ceiling_157,ceiling_154]=True
  close_item[ceiling_157,bathroom_cabinet_168]=True
  close_item[ceiling_157,faucet_172]=True
  close_item[ceiling_157,wall_151]=True
  close_item[ceiling_157,wall_152]=True
  close_item[ceiling_157,wall_153]=True
  close_item[ceiling_157,drawing_186]=True
  close_item[ceiling_157,ceiling_156]=True
  inside[tablelamp_317,home_office_248]=True
  on[nightstand_255,floor_341]=True
  on[plate_1005,kitchen_counter_1000]=True
  close_item[nightstand_72,doorjamb_228]=True
  close_item[nightstand_72,floor_5]=True
  close_item[nightstand_72,powersocket_197]=True
  close_item[nightstand_72,door_229]=True
  close_item[nightstand_72,orchid_136]=True
  close_item[nightstand_72,floor_8]=True
  close_item[nightstand_72,drawing_138]=True
  close_item[nightstand_72,couch_71]=True
  close_item[nightstand_72,floor_235]=True
  close_item[nightstand_72,floor_234]=True
  close_item[nightstand_72,wall_243]=True
  close_item[nightstand_72,wall_23]=True
  close_item[nightstand_72,wall_30]=True
  facing_item[ceilinglamp_34,drawing_139]=True
  facing_item[ceilinglamp_34,drawing_140]=True
  facing_item[ceilinglamp_34,drawing_141]=True
  facing_item[ceilinglamp_34,drawing_142]=True
  close_item[closetdrawer_267,dresser_258]=True
  close_item[closetdrawer_267,hanger_259]=True
  close_item[closetdrawer_267,hanger_260]=True
  close_item[closetdrawer_267,hanger_261]=True
  close_item[closetdrawer_267,hanger_262]=True
  close_item[closetdrawer_267,hanger_263]=True
  close_item[closetdrawer_267,hanger_264]=True
  close_item[closetdrawer_267,hanger_265]=True
  close_item[closetdrawer_267,closetdrawer_266]=True
  close_item[closetdrawer_267,closetdrawer_268]=True
  close_item[closetdrawer_267,closetdrawer_269]=True
  close_item[closetdrawer_267,closetdrawer_270]=True
  close_item[closetdrawer_267,closetdrawer_271]=True
  close_item[closetdrawer_267,closetdrawer_272]=True
  close_item[closetdrawer_267,television_278]=True
  close_item[closetdrawer_267,curtain_284]=True
  close_item[closetdrawer_267,curtain_285]=True
  close_item[closetdrawer_267,walllamp_315]=True
  close_item[closetdrawer_267,wall_321]=True
  close_item[closetdrawer_267,wall_325]=True
  close_item[closetdrawer_267,floor_343]=True
  close_item[closetdrawer_267,floor_344]=True
  close_item[closetdrawer_267,window_348]=True
  close_item[closetdrawer_267,tvstand_252]=True
  inside[couch_71,dining_room_1]=True
  inside[food_food_2016,cupboard_65]=True
  inside[food_food_2016,dining_room_1]=True
  inside[hanger_265,home_office_248]=True
  inside[hanger_265,dresser_258]=True
  facing_item[ceiling_332,drawing_283]=True
  facing_item[ceiling_332,television_278]=True
  facing_item[mat_185,drawing_186]=True
  inside[juice_2026,dining_room_1]=True
  inside[juice_2026,sink_67]=True
  close_item[floor_236,desk_192]=True
  close_item[floor_236,wall_322]=True
  close_item[floor_236,filing_cabinet_195]=True
  close_item[floor_236,mat_230]=True
  close_item[floor_236,floor_234]=True
  close_item[floor_236,floor_235]=True
  close_item[floor_236,photoframe_204]=True
  close_item[floor_236,floor_237]=True
  close_item[floor_236,floor_338]=True
  close_item[floor_236,wall_243]=True
  close_item[floor_236,wall_245]=True
  close_item[floor_236,wall_246]=True
  close_item[floor_236,light_280]=True
  close_item[floor_236,bookshelf_250]=True
  close_item[floor_236,door_347]=True
  close_item[floor_236,bookshelf_190]=True
  close_item[floor_236,chair_191]=True
  close_item[desk_251,wall_322]=True
  close_item[desk_251,keyboard_2057]=True
  close_item[desk_251,computer_273]=True
  close_item[desk_251,cpuscreen_274]=True
  close_item[desk_251,keyboard_275]=True
  close_item[desk_251,mousepad_276]=True
  close_item[desk_251,mouse_277]=True
  close_item[desk_251,floor_339]=True
  close_item[desk_251,walllamp_311]=True
  close_item[desk_251,walllamp_312]=True
  close_item[desk_251,floor_338]=True
  close_item[desk_251,cup_2010]=True
  close_item[desk_251,chair_254]=True
  close_item[desk_251,wall_319]=True
  inside[floor_336,home_office_248]=True
  close_item[form_2048,filing_cabinet_195]=True
  close_item[ceiling_20,ceilinglamp_35]=True
  close_item[ceiling_20,doorjamb_228]=True
  close_item[ceiling_20,wallshelf_74]=True
  close_item[ceiling_20,wallshelf_75]=True
  close_item[ceiling_20,drawing_138]=True
  close_item[ceiling_20,drawing_140]=True
  close_item[ceiling_20,curtain_143]=True
  close_item[ceiling_20,curtain_144]=True
  close_item[ceiling_20,ceiling_16]=True
  close_item[ceiling_20,ceiling_18]=True
  close_item[ceiling_20,ceiling_239]=True
  close_item[ceiling_20,wall_243]=True
  close_item[ceiling_20,wall_30]=True
  on[form_2015,bookshelf_190]=True
  on[check_2003,couch_256]=True
  close_item[clothes_dress_2007,couch_257]=True
  inside[floor_3,dining_room_1]=True
  inside[newspaper_2051,home_office_248]=True
  close_item[thread_2012,filing_cabinet_195]=True
  on[mouse_277,desk_251]=True
  on[mouse_277,mousepad_276]=True
  inside[wall_320,home_office_248]=True
  on[pillow_232,bed_194]=True
  close_item[couch_257,pillow_289]=True
  close_item[couch_257,pillow_290]=True
  close_item[couch_257,clothes_underwear_2049]=True
  close_item[couch_257,wall_324]=True
  close_item[couch_257,newspaper_2051]=True
  close_item[couch_257,ceiling_332]=True
  close_item[couch_257,walllamp_314]=True
  close_item[couch_257,floor_341]=True
  close_item[couch_257,floor_342]=True
  close_item[couch_257,clothes_dress_2007]=True
  close_item[couch_257,hanger_2014]=True
  close_item[couch_257,table_249]=True
  close_item[couch_257,orchid_282]=True
  close_item[couch_257,walllamp_316]=True
  close_item[couch_257,tablelamp_317]=True
  close_item[couch_257,wall_318]=True
  close_item[couch_257,nightstand_255]=True
  close_item[television_278,wall_321]=True
  close_item[television_278,dresser_258]=True
  close_item[television_278,wall_325]=True
  close_item[television_278,closetdrawer_267]=True
  close_item[television_278,closetdrawer_268]=True
  close_item[television_278,ceiling_333]=True
  close_item[television_278,closetdrawer_271]=True
  close_item[television_278,floor_339]=True
  close_item[television_278,tvstand_252]=True
  close_item[television_278,window_348]=True
  close_item[television_278,floor_340]=True
  close_item[television_278,floor_343]=True
  close_item[television_278,floor_344]=True
  close_item[television_278,table_249]=True
  close_item[television_278,walllamp_315]=True
  close_item[television_278,curtain_284]=True
  close_item[television_278,curtain_285]=True
  inside[curtain_284,home_office_248]=True
  inside[curtain_284,curtain_285]=True
  inside[food_butter_2035,dining_room_1]=True
  inside[food_butter_2035,microwave_86]=True
  close_item[orchid_282,couch_257]=True
  close_item[orchid_282,wall_321]=True
  close_item[orchid_282,wall_324]=True
  close_item[orchid_282,floor_340]=True
  close_item[orchid_282,floor_341]=True
  close_item[orchid_282,floor_342]=True
  close_item[orchid_282,floor_343]=True
  close_item[orchid_282,table_249]=True
  close_item[orchid_282,tvstand_252]=True
  close_item[orchid_282,curtain_286]=True
  inside[coffe_maker_84,dining_room_1]=True
  close_item[ceiling_326,wall_323]=True
  close_item[ceiling_326,light_196]=True
  close_item[ceiling_326,photoframe_294]=True
  close_item[ceiling_326,ceiling_327]=True
  close_item[ceiling_326,ceiling_331]=True
  close_item[ceiling_326,ceilinglamp_310]=True
  close_item[ceiling_326,walllamp_313]=True
  close_item[ceiling_326,walllamp_314]=True
  close_item[ceiling_326,drawing_283]=True
  close_item[ceiling_326,bookshelf_253]=True
  inside[ceiling_12,dining_room_1]=True
  inside[napkin_2019,cupboard_64]=True
  inside[napkin_2019,dining_room_1]=True
  inside[ground_coffee_2060,dining_room_1]=True
  inside[ground_coffee_2060,coffe_maker_84]=True
  close_item[ceiling_330,couch_256]=True
  close_item[ceiling_330,ceiling_327]=True
  close_item[ceiling_330,ceiling_329]=True
  close_item[ceiling_330,ceiling_331]=True
  close_item[ceiling_330,ceiling_333]=True
  close_item[ceiling_330,ceilinglamp_310]=True
  inside[doorjamb_32,dining_room_1]=True
  inside[ceiling_329,home_office_248]=True
  facing_item[mat_135,drawing_139]=True
  facing_item[mat_135,drawing_140]=True
  facing_item[mat_135,drawing_141]=True
  facing_item[mat_135,drawing_142]=True
  inside[tvstand_252,home_office_248]=True
  on[closetdrawer_266,closetdrawer_269]=True
  close_item[chair_59,ceilinglamp_34]=True
  close_item[chair_59,floor_2]=True
  close_item[chair_59,floor_4]=True
  close_item[chair_59,floor_5]=True
  close_item[chair_59,floor_3]=True
  close_item[chair_59,floor_7]=True
  close_item[chair_59,floor_6]=True
  close_item[chair_59,wall_22]=True
  close_item[chair_59,wall_30]=True
  close_item[chair_59,chair_60]=True
  close_item[chair_59,chair_61]=True
  close_item[chair_59,chair_62]=True
  close_item[chair_59,table_63]=True
  facing_item[ceiling_14,drawing_139]=True
  facing_item[ceiling_14,drawing_140]=True
  facing_item[ceiling_14,drawing_141]=True
  facing_item[ceiling_14,drawing_142]=True
  on[closetdrawer_270,closetdrawer_272]=True
  facing_item[bathroom_counter_171,drawing_186]=True
  close_item[stovefan_79,cupboard_64]=True
  close_item[stovefan_79,pot_97]=True
  close_item[stovefan_79,pot_98]=True
  close_item[stovefan_79,cupboard_65]=True
  close_item[stovefan_79,walllamp_36]=True
  close_item[stovefan_79,kitchen_counter_69]=True
  close_item[stovefan_79,kitchen_counter_66]=True
  close_item[stovefan_79,ceiling_12]=True
  close_item[stovefan_79,toaster_76]=True
  close_item[stovefan_79,ceiling_13]=True
  close_item[stovefan_79,oven_82]=True
  close_item[stovefan_79,tray_83]=True
  close_item[stovefan_79,ceiling_19]=True
  close_item[stovefan_79,wall_21]=True
  close_item[stovefan_79,wall_24]=True
  close_item[stovefan_79,wall_25]=True
  close_item[stovefan_79,wall_26]=True
  close_item[stovefan_79,knifeblock_92]=True
  close_item[stovefan_79,wall_29]=True
  close_item[coffe_maker_84,cupboard_64]=True
  close_item[coffe_maker_84,kitchen_counter_69]=True
  close_item[coffe_maker_84,kitchen_counter_70]=True
  close_item[coffe_maker_84,floor_10]=True
  close_item[coffe_maker_84,ground_coffee_2060]=True
  close_item[coffe_maker_84,dishwasher_81]=True
  close_item[coffe_maker_84,ceiling_19]=True
  close_item[coffe_maker_84,wall_25]=True
  close_item[coffe_maker_84,wall_26]=True
  close_item[coffe_maker_84,wall_29]=True
  inside[sink_67,dining_room_1]=True
  inside[sink_67,kitchen_counter_66]=True
  inside[mouse_277,home_office_248]=True
  inside[check_2002,home_office_248]=True
  inside[door_31,dining_room_1]=True
  close_item[wall_321,dresser_258]=True
  close_item[wall_321,hanger_259]=True
  close_item[wall_321,hanger_260]=True
  close_item[wall_321,hanger_261]=True
  close_item[wall_321,closetdrawer_267]=True
  close_item[wall_321,closetdrawer_268]=True
  close_item[wall_321,closetdrawer_271]=True
  close_item[wall_321,television_278]=True
  close_item[wall_321,orchid_282]=True
  close_item[wall_321,curtain_284]=True
  close_item[wall_321,curtain_285]=True
  close_item[wall_321,curtain_286]=True
  close_item[wall_321,walllamp_315]=True
  close_item[wall_321,walllamp_316]=True
  close_item[wall_321,wall_324]=True
  close_item[wall_321,wall_325]=True
  close_item[wall_321,ceiling_333]=True
  close_item[wall_321,floor_343]=True
  close_item[wall_321,window_348]=True
  close_item[wall_321,table_249]=True
  close_item[wall_321,tvstand_252]=True
  close_item[floor_341,couch_256]=True
  close_item[floor_341,pillow_288]=True
  close_item[floor_341,pillow_289]=True
  close_item[floor_341,couch_257]=True
  close_item[floor_341,pillow_287]=True
  close_item[floor_341,wall_324]=True
  close_item[floor_341,wall_323]=True
  close_item[floor_341,orchid_282]=True
  close_item[floor_341,floor_335]=True
  close_item[floor_341,floor_336]=True
  close_item[floor_341,floor_340]=True
  close_item[floor_341,floor_342]=True
  close_item[floor_341,table_249]=True
  close_item[floor_341,walllamp_314]=True
  close_item[floor_341,drawing_283]=True
  close_item[floor_341,tablelamp_317]=True
  close_item[floor_341,wall_318]=True
  close_item[floor_341,nightstand_255]=True
  on[pencil_2039,table_249]=True
  close_item[doorjamb_346,dresser_258]=True
  close_item[doorjamb_346,hanger_259]=True
  close_item[doorjamb_346,hanger_260]=True
  close_item[doorjamb_346,wall_325]=True
  close_item[doorjamb_346,hanger_262]=True
  close_item[doorjamb_346,hanger_263]=True
  close_item[doorjamb_346,hanger_264]=True
  close_item[doorjamb_346,hanger_265]=True
  close_item[doorjamb_346,closetdrawer_266]=True
  close_item[doorjamb_346,hanger_261]=True
  close_item[doorjamb_346,closetdrawer_269]=True
  close_item[doorjamb_346,closetdrawer_270]=True
  close_item[doorjamb_346,ceiling_334]=True
  close_item[doorjamb_346,closetdrawer_272]=True
  close_item[doorjamb_346,floor_344]=True
  close_item[doorjamb_346,wall_319]=True
  inside[floor_235,bedroom_189]=True
  facing_item[ceiling_326,drawing_283]=True
  inside[ceiling_15,dining_room_1]=True
  inside[after_shave_2063,dining_room_1]=True
  inside[after_shave_2063,sink_67]=True
  close_item[photoframe_133,floor_161]=True
  close_item[photoframe_133,floor_6]=True
  close_item[photoframe_133,couch_71]=True
  close_item[photoframe_133,shower_167]=True
  close_item[photoframe_133,nightstand_73]=True
  close_item[photoframe_133,shower_169]=True
  close_item[photoframe_133,drawing_142]=True
  close_item[photoframe_133,freezer_80]=True
  close_item[photoframe_133,wall_22]=True
  close_item[photoframe_133,wall_153]=True
  close_item[drawing_138,couch_71]=True
  close_item[drawing_138,orchid_136]=True
  close_item[drawing_138,nightstand_72]=True
  close_item[drawing_138,drawing_139]=True
  close_item[drawing_138,drawing_140]=True
  close_item[drawing_138,drawing_141]=True
  close_item[drawing_138,ceiling_239]=True
  close_item[drawing_138,ceiling_16]=True
  close_item[drawing_138,wall_243]=True
  close_item[drawing_138,ceiling_20]=True
  close_item[drawing_138,wall_22]=True
  close_item[drawing_138,wall_23]=True
  close_item[drawing_138,wall_30]=True
  close_item[curtain_144,window_33]=True
  close_item[curtain_144,floor_7]=True
  close_item[curtain_144,wallshelf_74]=True
  close_item[curtain_144,wallshelf_75]=True
  close_item[curtain_144,curtain_143]=True
  close_item[curtain_144,curtain_145]=True
  close_item[curtain_144,ceiling_18]=True
  close_item[curtain_144,ceiling_20]=True
  close_item[curtain_144,wall_27]=True
  close_item[curtain_144,wall_30]=True
  inside[hanger_260,home_office_248]=True
  inside[hanger_260,dresser_258]=True
  close_item[oven_82,cupboard_64]=True
  close_item[oven_82,pot_97]=True
  close_item[oven_82,pot_98]=True
  close_item[oven_82,kitchen_counter_66]=True
  close_item[oven_82,walllamp_36]=True
  close_item[oven_82,kitchen_counter_69]=True
  close_item[oven_82,cupboard_65]=True
  close_item[oven_82,floor_9]=True
  close_item[oven_82,floor_11]=True
  close_item[oven_82,toaster_76]=True
  close_item[oven_82,ceiling_12]=True
  close_item[oven_82,stovefan_79]=True
  close_item[oven_82,tray_83]=True
  close_item[oven_82,wall_21]=True
  close_item[oven_82,wall_24]=True
  close_item[oven_82,wall_25]=True
  close_item[oven_82,wall_26]=True
  close_item[oven_82,knifeblock_92]=True
  close_item[oven_82,wall_29]=True
  close_item[pot_97,cupboard_64]=True
  close_item[pot_97,cupboard_65]=True
  close_item[pot_97,pot_98]=True
  close_item[pot_97,kitchen_counter_66]=True
  close_item[pot_97,walllamp_36]=True
  close_item[pot_97,kitchen_counter_69]=True
  close_item[pot_97,floor_11]=True
  close_item[pot_97,toaster_76]=True
  close_item[pot_97,ceiling_12]=True
  close_item[pot_97,stovefan_79]=True
  close_item[pot_97,dishwasher_81]=True
  close_item[pot_97,oven_82]=True
  close_item[pot_97,tray_83]=True
  close_item[pot_97,wall_21]=True
  close_item[pot_97,wall_24]=True
  close_item[pot_97,wall_25]=True
  close_item[pot_97,wall_26]=True
  close_item[pot_97,knifeblock_92]=True
  close_item[pot_97,wall_29]=True
  inside[chair_60,dining_room_1]=True
  on[closetdrawer_267,closetdrawer_268]=True
  close_item[tablelamp_317,couch_256]=True
  close_item[tablelamp_317,pillow_289]=True
  close_item[tablelamp_317,pillow_288]=True
  close_item[tablelamp_317,couch_257]=True
  close_item[tablelamp_317,wall_324]=True
  close_item[tablelamp_317,wall_323]=True
  close_item[tablelamp_317,ceiling_331]=True
  close_item[tablelamp_317,floor_341]=True
  close_item[tablelamp_317,floor_342]=True
  close_item[tablelamp_317,walllamp_314]=True
  close_item[tablelamp_317,drawing_283]=True
  close_item[tablelamp_317,wall_318]=True
  close_item[tablelamp_317,nightstand_255]=True
  inside[floor_8,dining_room_1]=True
  inside[detergent_2056,filing_cabinet_195]=True
  inside[detergent_2056,bedroom_189]=True
  on[clothes_hat_2028,couch_71]=True
  close_item[window_348,wall_321]=True
  close_item[window_348,dresser_258]=True
  close_item[window_348,hanger_259]=True
  close_item[window_348,hanger_260]=True
  close_item[window_348,wall_324]=True
  close_item[window_348,wall_325]=True
  close_item[window_348,closetdrawer_267]=True
  close_item[window_348,closetdrawer_268]=True
  close_item[window_348,ceiling_333]=True
  close_item[window_348,closetdrawer_271]=True
  close_item[window_348,floor_343]=True
  close_item[window_348,tvstand_252]=True
  close_item[window_348,walllamp_316]=True
  close_item[window_348,television_278]=True
  close_item[window_348,walllamp_315]=True
  close_item[window_348,curtain_284]=True
  close_item[window_348,curtain_285]=True
  close_item[window_348,curtain_286]=True
  inside[ceiling_18,dining_room_1]=True
  inside[shoes_2066,home_office_248]=True
  inside[shoes_2066,dresser_258]=True
  inside[doorjamb_228,bedroom_189]=True
  facing_item[ceiling_333,computer_273]=True
  facing_item[ceiling_333,television_278]=True
  facing_item[doorjamb_345,computer_273]=True
  facing_item[doorjamb_345,drawing_283]=True
  close_item[hanger_259,dresser_258]=True
  close_item[hanger_259,hanger_260]=True
  close_item[hanger_259,hanger_261]=True
  close_item[hanger_259,hanger_262]=True
  close_item[hanger_259,hanger_263]=True
  close_item[hanger_259,hanger_264]=True
  close_item[hanger_259,hanger_265]=True
  close_item[hanger_259,closetdrawer_266]=True
  close_item[hanger_259,closetdrawer_267]=True
  close_item[hanger_259,closetdrawer_268]=True
  close_item[hanger_259,closetdrawer_269]=True
  close_item[hanger_259,closetdrawer_270]=True
  close_item[hanger_259,curtain_284]=True
  close_item[hanger_259,curtain_285]=True
  close_item[hanger_259,walllamp_315]=True
  close_item[hanger_259,wall_321]=True
  close_item[hanger_259,wall_325]=True
  close_item[hanger_259,ceiling_333]=True
  close_item[hanger_259,ceiling_334]=True
  close_item[hanger_259,doorjamb_346]=True
  close_item[hanger_259,window_348]=True
  close_item[powersocket_197,nightstand_193]=True
  close_item[powersocket_197,doorjamb_228]=True
  close_item[powersocket_197,door_229]=True
  close_item[powersocket_197,floor_5]=True
  close_item[powersocket_197,mat_230]=True
  close_item[powersocket_197,nightstand_72]=True
  close_item[powersocket_197,orchid_136]=True
  close_item[powersocket_197,floor_234]=True
  close_item[powersocket_197,floor_235]=True
  close_item[powersocket_197,floor_8]=True
  close_item[powersocket_197,couch_71]=True
  close_item[powersocket_197,wall_243]=True
  close_item[powersocket_197,wall_23]=True
  close_item[powersocket_197,bookshelf_190]=True
  close_item[powersocket_197,wall_30]=True
  inside[floor_160,bathroom_149]=True
  facing_item[floor_7,drawing_138]=True
  facing_item[floor_7,drawing_139]=True
  facing_item[floor_7,drawing_140]=True
  inside[wall_27,dining_room_1]=True
  close_item[doorjamb_228,nightstand_193]=True
  close_item[doorjamb_228,powersocket_197]=True
  close_item[doorjamb_228,door_229]=True
  close_item[doorjamb_228,orchid_136]=True
  close_item[doorjamb_228,floor_8]=True
  close_item[doorjamb_228,floor_234]=True
  close_item[doorjamb_228,floor_235]=True
  close_item[doorjamb_228,nightstand_72]=True
  close_item[doorjamb_228,wallshelf_75]=True
  close_item[doorjamb_228,ceiling_239]=True
  close_item[doorjamb_228,wall_243]=True
  close_item[doorjamb_228,ceiling_20]=True
  close_item[doorjamb_228,wall_244]=True
  close_item[doorjamb_228,wall_23]=True
  close_item[doorjamb_228,bookshelf_190]=True
  close_item[doorjamb_228,wall_30]=True
  on[nightstand_72,floor_5]=True
  between[door_229,dining_room_1]=True
  between[door_229,bedroom_189]=True
  close_item[wall_243,orchid_136]=True
  close_item[wall_243,floor_8]=True
  close_item[wall_243,drawing_138]=True
  close_item[wall_243,drawing_140]=True
  close_item[wall_243,ceiling_20]=True
  close_item[wall_243,wall_23]=True
  close_item[wall_243,wall_30]=True
  close_item[wall_243,bookshelf_190]=True
  close_item[wall_243,chair_191]=True
  close_item[wall_243,nightstand_193]=True
  close_item[wall_243,bed_194]=True
  close_item[wall_243,powersocket_197]=True
  close_item[wall_243,nightstand_72]=True
  close_item[wall_243,photoframe_204]=True
  close_item[wall_243,doorjamb_228]=True
  close_item[wall_243,door_229]=True
  close_item[wall_243,mat_230]=True
  close_item[wall_243,pillow_231]=True
  close_item[wall_243,ceilinglamp_233]=True
  close_item[wall_243,floor_234]=True
  close_item[wall_243,floor_235]=True
  close_item[wall_243,floor_236]=True
  close_item[wall_243,floor_238]=True
  close_item[wall_243,ceiling_239]=True
  close_item[wall_243,ceiling_240]=True
  close_item[wall_243,ceiling_242]=True
  close_item[wall_243,wall_244]=True
  close_item[wall_243,wall_245]=True
  inside_char[char,bedroom_189]=True
  on[wall_24,kitchen_counter_66]=True
  facing_item[bathroom_cabinet_168,drawing_186]=True
  close_item[wall_151,floor_160]=True
  close_item[wall_151,floor_162]=True
  close_item[wall_151,walllamp_163]=True
  close_item[wall_151,ceilinglamp_164]=True
  close_item[wall_151,bathroom_cabinet_168]=True
  close_item[wall_151,bathroom_counter_171]=True
  close_item[wall_151,faucet_172]=True
  close_item[wall_151,sink_173]=True
  close_item[wall_151,wall_150]=True
  close_item[wall_151,wall_152]=True
  close_item[wall_151,mat_185]=True
  close_item[wall_151,ceiling_154]=True
  close_item[wall_151,ceiling_155]=True
  close_item[wall_151,ceiling_157]=True
  close_item[wall_151,floor_158]=True
  close_item[wall_151,floor_159]=True
  inside[filing_cabinet_195,bedroom_189]=True
  close_item[food_peanut_butter_2022,cupboard_65]=True
  close_item[ceiling_156,ceilinglamp_164]=True
  close_item[ceiling_156,shower_167]=True
  close_item[ceiling_156,shower_169]=True
  close_item[ceiling_156,curtain_170]=True
  close_item[ceiling_156,ceiling_17]=True
  close_item[ceiling_156,light_146]=True
  close_item[ceiling_156,wall_150]=True
  close_item[ceiling_156,wall_22]=True
  close_item[ceiling_156,wall_152]=True
  close_item[ceiling_156,wall_153]=True
  close_item[ceiling_156,drawing_186]=True
  close_item[ceiling_156,ceiling_155]=True
  close_item[ceiling_156,ceiling_157]=True
  close_item[homework_2027,filing_cabinet_195]=True
  inside[pillow_231,bedroom_189]=True
  close_item[dvd_player_2047,table_249]=True
  close_item[closetdrawer_270,dresser_258]=True
  close_item[closetdrawer_270,hanger_259]=True
  close_item[closetdrawer_270,hanger_260]=True
  close_item[closetdrawer_270,wall_325]=True
  close_item[closetdrawer_270,hanger_262]=True
  close_item[closetdrawer_270,hanger_263]=True
  close_item[closetdrawer_270,hanger_261]=True
  close_item[closetdrawer_270,hanger_265]=True
  close_item[closetdrawer_270,closetdrawer_266]=True
  close_item[closetdrawer_270,closetdrawer_267]=True
  close_item[closetdrawer_270,closetdrawer_268]=True
  close_item[closetdrawer_270,closetdrawer_269]=True
  close_item[closetdrawer_270,hanger_264]=True
  close_item[closetdrawer_270,closetdrawer_271]=True
  close_item[closetdrawer_270,closetdrawer_272]=True
  close_item[closetdrawer_270,floor_344]=True
  close_item[closetdrawer_270,doorjamb_346]=True
  close_item[closetdrawer_270,walllamp_315]=True
  inside[floor_159,bathroom_149]=True
  on[ceiling_17,wall_22]=True
  close_item[photoframe_204,desk_192]=True
  close_item[photoframe_204,mat_230]=True
  close_item[photoframe_204,floor_234]=True
  close_item[photoframe_204,floor_235]=True
  close_item[photoframe_204,floor_236]=True
  close_item[photoframe_204,ceiling_239]=True
  close_item[photoframe_204,ceiling_240]=True
  close_item[photoframe_204,wall_243]=True
  close_item[photoframe_204,wall_245]=True
  close_item[photoframe_204,bookshelf_190]=True
  close_item[photoframe_204,chair_191]=True
  close_item[wall_318,couch_256]=True
  close_item[wall_318,pillow_289]=True
  close_item[wall_318,couch_257]=True
  close_item[wall_318,wall_323]=True
  close_item[wall_318,wall_324]=True
  close_item[wall_318,ceiling_331]=True
  close_item[wall_318,floor_341]=True
  close_item[wall_318,walllamp_313]=True
  close_item[wall_318,walllamp_314]=True
  close_item[wall_318,drawing_283]=True
  close_item[wall_318,tablelamp_317]=True
  close_item[wall_318,nightstand_255]=True
  on[sponge_2040,bathroom_counter_171]=True
  inside[curtain_143,curtain_144]=True
  inside[curtain_143,dining_room_1]=True
  close_item[floor_6,floor_161]=True
  close_item[floor_6,floor_2]=True
  close_item[floor_6,floor_3]=True
  close_item[floor_6,photoframe_133]=True
  close_item[floor_6,toilet_166]=True
  close_item[floor_6,couch_71]=True
  close_item[floor_6,floor_5]=True
  close_item[floor_6,nightstand_73]=True
  close_item[floor_6,shower_169]=True
  close_item[floor_6,mat_135]=True
  close_item[floor_6,shower_167]=True
  close_item[floor_6,freezer_80]=True
  close_item[floor_6,light_146]=True
  close_item[floor_6,powersocket_147]=True
  close_item[floor_6,wall_22]=True
  close_item[floor_6,wall_153]=True
  close_item[floor_6,chair_59]=True
  close_item[floor_6,door_31]=True
  close_item[check_2054,filing_cabinet_195]=True
  close_item[door_31,doorjamb_32]=True
  close_item[door_31,floor_160]=True
  close_item[door_31,floor_2]=True
  close_item[door_31,floor_3]=True
  close_item[door_31,floor_161]=True
  close_item[door_31,toilet_166]=True
  close_item[door_31,mat_135]=True
  close_item[door_31,shower_167]=True
  close_item[door_31,floor_9]=True
  close_item[door_31,floor_6]=True
  close_item[door_31,freezer_80]=True
  close_item[door_31,light_146]=True
  close_item[door_31,powersocket_147]=True
  close_item[door_31,wall_21]=True
  close_item[door_31,wall_150]=True
  close_item[door_31,wall_22]=True
  close_item[door_31,wall_153]=True
  close_item[door_31,light_187]=True
  close_item[door_31,wall_28]=True
  inside[door_347,home_office_248]=True
  on[clothes_scarf_2004,couch_71]=True
  on[food_food_2033,plate_1005]=True
  close_item[couch_256,pillow_287]=True
  close_item[couch_256,pillow_288]=True
  close_item[couch_256,pillow_289]=True
  close_item[couch_256,ceilinglamp_310]=True
  close_item[couch_256,walllamp_314]=True
  close_item[couch_256,tablelamp_317]=True
  close_item[couch_256,wall_318]=True
  close_item[couch_256,wall_323]=True
  close_item[couch_256,wall_324]=True
  close_item[couch_256,ceiling_330]=True
  close_item[couch_256,ceiling_331]=True
  close_item[couch_256,floor_335]=True
  close_item[couch_256,floor_336]=True
  close_item[couch_256,floor_337]=True
  close_item[couch_256,check_2003]=True
  close_item[couch_256,floor_340]=True
  close_item[couch_256,floor_341]=True
  close_item[couch_256,floor_342]=True
  close_item[couch_256,floor_343]=True
  close_item[couch_256,tray_2021]=True
  close_item[couch_256,clothes_shirt_2038]=True
  close_item[couch_256,chair_254]=True
  close_item[couch_256,nightstand_255]=True
  close_item[bed_194,nightstand_193]=True
  close_item[bed_194,mat_230]=True
  close_item[bed_194,pillow_231]=True
  close_item[bed_194,pillow_232]=True
  close_item[bed_194,floor_234]=True
  close_item[bed_194,floor_235]=True
  close_item[bed_194,floor_237]=True
  close_item[bed_194,floor_238]=True
  close_item[bed_194,sheets_2032]=True
  close_item[bed_194,wall_243]=True
  close_item[bed_194,wall_244]=True
  close_item[bed_194,wall_246]=True
  inside[orchid_136,dining_room_1]=True
  inside[bookmark_2046,filing_cabinet_195]=True
  inside[bookmark_2046,bedroom_189]=True
  inside[light_146,dining_room_1]=True
  close_item[ceiling_242,ceilinglamp_233]=True
  close_item[ceiling_242,ceiling_239]=True
  close_item[ceiling_242,ceiling_241]=True
  close_item[ceiling_242,wall_243]=True
  close_item[ceiling_242,wall_244]=True
  close_item[ceiling_242,wall_246]=True
  close_item[floor_7,floor_4]=True
  close_item[floor_7,floor_8]=True
  close_item[floor_7,chair_59]=True
  close_item[floor_7,floor_10]=True
  close_item[floor_7,curtain_143]=True
  close_item[floor_7,curtain_144]=True
  close_item[floor_7,curtain_145]=True
  close_item[floor_7,wall_29]=True
  close_item[floor_7,wall_30]=True
  close_item[floor_7,wall_27]=True
  close_item[floor_7,chair_60]=True
  close_item[floor_7,chair_61]=True
  close_item[floor_7,chair_62]=True
  close_item[floor_7,table_63]=True
  close_item[band_aids_2055,bathroom_counter_171]=True
  facing_item[ceiling_330,computer_273]=True
  facing_item[ceiling_330,drawing_283]=True
  inside[floor_340,home_office_248]=True
  close_item[shoe_rack_2013,mat_230]=True
  close_item[food_carrot_2018,plate_1004]=True
  close_item[orchid_136,doorjamb_228]=True
  close_item[orchid_136,door_229]=True
  close_item[orchid_136,floor_5]=True
  close_item[orchid_136,powersocket_197]=True
  close_item[orchid_136,nightstand_72]=True
  close_item[orchid_136,floor_8]=True
  close_item[orchid_136,drawing_138]=True
  close_item[orchid_136,couch_71]=True
  close_item[orchid_136,floor_235]=True
  close_item[orchid_136,floor_234]=True
  close_item[orchid_136,wall_243]=True
  close_item[orchid_136,wall_23]=True
  close_item[orchid_136,wall_30]=True
  inside[pillow_288,home_office_248]=True
  inside[ceiling_155,bathroom_149]=True
  close_item[closetdrawer_269,dresser_258]=True
  close_item[closetdrawer_269,hanger_259]=True
  close_item[closetdrawer_269,hanger_260]=True
  close_item[closetdrawer_269,wall_325]=True
  close_item[closetdrawer_269,hanger_262]=True
  close_item[closetdrawer_269,hanger_263]=True
  close_item[closetdrawer_269,hanger_261]=True
  close_item[closetdrawer_269,hanger_265]=True
  close_item[closetdrawer_269,closetdrawer_266]=True
  close_item[closetdrawer_269,closetdrawer_267]=True
  close_item[closetdrawer_269,closetdrawer_268]=True
  close_item[closetdrawer_269,hanger_264]=True
  close_item[closetdrawer_269,closetdrawer_270]=True
  close_item[closetdrawer_269,closetdrawer_271]=True
  close_item[closetdrawer_269,closetdrawer_272]=True
  close_item[closetdrawer_269,floor_344]=True
  close_item[closetdrawer_269,doorjamb_346]=True
  close_item[closetdrawer_269,walllamp_315]=True
  facing_item[wall_150,drawing_186]=True
  inside[plate_1005,dishwasher_1002]=True
  inside[plate_1005,bedroom_189]=True
  facing_item[floor_4,drawing_138]=True
  facing_item[floor_4,drawing_139]=True
  facing_item[floor_4,drawing_140]=True
  facing_item[floor_4,drawing_141]=True
  facing_item[floor_4,drawing_142]=True
  close_item[walllamp_315,dresser_258]=True
  close_item[walllamp_315,hanger_259]=True
  close_item[walllamp_315,hanger_260]=True
  close_item[walllamp_315,hanger_261]=True
  close_item[walllamp_315,hanger_262]=True
  close_item[walllamp_315,hanger_263]=True
  close_item[walllamp_315,hanger_265]=True
  close_item[walllamp_315,closetdrawer_266]=True
  close_item[walllamp_315,closetdrawer_267]=True
  close_item[walllamp_315,closetdrawer_268]=True
  close_item[walllamp_315,closetdrawer_269]=True
  close_item[walllamp_315,closetdrawer_270]=True
  close_item[walllamp_315,closetdrawer_271]=True
  close_item[walllamp_315,closetdrawer_272]=True
  close_item[walllamp_315,television_278]=True
  close_item[walllamp_315,curtain_284]=True
  close_item[walllamp_315,curtain_285]=True
  close_item[walllamp_315,wall_321]=True
  close_item[walllamp_315,wall_325]=True
  close_item[walllamp_315,ceiling_333]=True
  close_item[walllamp_315,ceiling_334]=True
  close_item[walllamp_315,floor_344]=True
  close_item[walllamp_315,window_348]=True
  close_item[walllamp_315,tvstand_252]=True
  on[bookmark_2053,desk_192]=True
  close_item[wall_320,wall_322]=True
  close_item[wall_320,filing_cabinet_195]=True
  close_item[wall_320,light_196]=True
  close_item[wall_320,wall_323]=True
  close_item[wall_320,mat_281]=True
  close_item[wall_320,ceiling_327]=True
  close_item[wall_320,photoframe_294]=True
  close_item[wall_320,floor_237]=True
  close_item[wall_320,floor_337]=True
  close_item[wall_320,ceiling_241]=True
  close_item[wall_320,wall_245]=True
  close_item[wall_320,wall_246]=True
  close_item[wall_320,powersocket_279]=True
  close_item[wall_320,light_280]=True
  close_item[wall_320,doorjamb_345]=True
  close_item[wall_320,bookshelf_250]=True
  close_item[wall_320,door_347]=True
  close_item[wall_320,bookshelf_253]=True
  inside[drawing_139,dining_room_1]=True
  on[table_249,floor_343]=True
  facing_item[wall_28,drawing_139]=True
  facing_item[wall_28,drawing_141]=True
  facing_item[wall_28,drawing_142]=True
  close_item[bookshelf_253,wall_320]=True
  close_item[bookshelf_253,wall_323]=True
  close_item[bookshelf_253,light_196]=True
  close_item[bookshelf_253,photoframe_294]=True
  close_item[bookshelf_253,ceiling_326]=True
  close_item[bookshelf_253,doorjamb_345]=True
  close_item[bookshelf_253,mat_281]=True
  close_item[bookshelf_253,ceiling_327]=True
  close_item[bookshelf_253,floor_237]=True
  close_item[bookshelf_253,floor_335]=True
  close_item[bookshelf_253,floor_336]=True
  close_item[bookshelf_253,floor_337]=True
  close_item[bookshelf_253,check_2002]=True
  close_item[bookshelf_253,wall_246]=True
  close_item[bookshelf_253,powersocket_279]=True
  close_item[bookshelf_253,walllamp_313]=True
  close_item[bookshelf_253,door_347]=True
  close_item[floor_2,doorjamb_32]=True
  close_item[floor_2,floor_160]=True
  close_item[floor_2,floor_3]=True
  close_item[floor_2,floor_4]=True
  close_item[floor_2,toilet_166]=True
  close_item[floor_2,mat_135]=True
  close_item[floor_2,floor_6]=True
  close_item[floor_2,floor_9]=True
  close_item[floor_2,chair_59]=True
  close_item[floor_2,shower_167]=True
  close_item[floor_2,freezer_80]=True
  close_item[floor_2,light_146]=True
  close_item[floor_2,powersocket_147]=True
  close_item[floor_2,wall_21]=True
  close_item[floor_2,wall_22]=True
  close_item[floor_2,wall_150]=True
  close_item[floor_2,light_187]=True
  close_item[floor_2,wall_28]=True
  close_item[floor_2,chair_61]=True
  close_item[floor_2,door_31]=True
  close_item[floor_340,couch_256]=True
  close_item[floor_340,pillow_288]=True
  close_item[floor_340,table_249]=True
  close_item[floor_340,floor_337]=True
  close_item[floor_340,floor_339]=True
  close_item[floor_340,floor_341]=True
  close_item[floor_340,television_278]=True
  close_item[floor_340,floor_343]=True
  close_item[floor_340,mat_281]=True
  close_item[floor_340,orchid_282]=True
  close_item[floor_340,tvstand_252]=True
  close_item[floor_340,chair_254]=True
  close_item[floor_340,pillow_287]=True
  inside[shoe_rack_2013,bedroom_189]=True
  close_item[coffee_filter_2050,kitchen_counter_66]=True
  inside[wall_323,home_office_248]=True
  facing_item[ceiling_18,drawing_138]=True
  facing_item[ceiling_18,drawing_139]=True
  facing_item[ceiling_18,drawing_140]=True
  facing_item[photoframe_133,drawing_141]=True
  facing_item[photoframe_133,drawing_142]=True
  on[tray_2021,couch_256]=True
  facing_item[walllamp_316,television_278]=True
  inside[phone_148,dining_room_1]=True
  close_item[filing_cabinet_195,form_2048]=True
  close_item[filing_cabinet_195,clothes_socks_2052]=True
  close_item[filing_cabinet_195,check_2054]=True
  close_item[filing_cabinet_195,detergent_2056]=True
  close_item[filing_cabinet_195,toothbrush_holder_2059]=True
  close_item[filing_cabinet_195,powersocket_279]=True
  close_item[filing_cabinet_195,light_280]=True
  close_item[filing_cabinet_195,mat_281]=True
  close_item[filing_cabinet_195,wall_320]=True
  close_item[filing_cabinet_195,desk_192]=True
  close_item[filing_cabinet_195,wall_322]=True
  close_item[filing_cabinet_195,light_196]=True
  close_item[filing_cabinet_195,floor_337]=True
  close_item[filing_cabinet_195,floor_338]=True
  close_item[filing_cabinet_195,oven_mitts_2005]=True
  close_item[filing_cabinet_195,needle_2009]=True
  close_item[filing_cabinet_195,doorjamb_345]=True
  close_item[filing_cabinet_195,cd_2011]=True
  close_item[filing_cabinet_195,thread_2012]=True
  close_item[filing_cabinet_195,door_347]=True
  close_item[filing_cabinet_195,homework_2027]=True
  close_item[filing_cabinet_195,floor_236]=True
  close_item[filing_cabinet_195,floor_237]=True
  close_item[filing_cabinet_195,wall_245]=True
  close_item[filing_cabinet_195,wall_246]=True
  close_item[filing_cabinet_195,detergent_2041]=True
  close_item[filing_cabinet_195,bookshelf_250]=True
  close_item[filing_cabinet_195,bookmark_2046]=True
  inside[closetdrawer_271,home_office_248]=True
  inside[closetdrawer_271,dresser_258]=True
  inside[food_peanut_butter_2022,cupboard_65]=True
  inside[food_peanut_butter_2022,dining_room_1]=True
  inside[dishwasher_81,dining_room_1]=True
  on[closetdrawer_268,closetdrawer_271]=True
  facing_item[shower_169,drawing_186]=True
  inside[food_orange_2042,freezer_80]=True
  inside[food_orange_2042,dining_room_1]=True
  on[coffe_maker_84,kitchen_counter_69]=True
  inside[detergent_2006,bathroom_cabinet_168]=True
  inside[detergent_2006,bathroom_149]=True
  facing_item[table_63,drawing_138]=True
  facing_item[table_63,drawing_139]=True
  facing_item[table_63,drawing_140]=True
  facing_item[table_63,drawing_141]=True
  facing_item[table_63,drawing_142]=True
  inside[ceiling_19,dining_room_1]=True
  inside[walllamp_316,home_office_248]=True
  inside[wooden_spoon_2067,dining_room_1]=True
  close_item[curtain_143,window_33]=True
  close_item[curtain_143,floor_7]=True
  close_item[curtain_143,wallshelf_74]=True
  close_item[curtain_143,wallshelf_75]=True
  close_item[curtain_143,curtain_144]=True
  close_item[curtain_143,curtain_145]=True
  close_item[curtain_143,ceiling_18]=True
  close_item[curtain_143,ceiling_20]=True
  close_item[curtain_143,wall_27]=True
  close_item[curtain_143,wall_30]=True
  close_item[hanger_2014,couch_257]=True
  close_item[phone_148,doorjamb_32]=True
  close_item[phone_148,cupboard_65]=True
  close_item[phone_148,kitchen_counter_66]=True
  close_item[phone_148,floor_9]=True
  close_item[phone_148,ceiling_155]=True
  close_item[phone_148,ceiling_13]=True
  close_item[phone_148,ceiling_14]=True
  close_item[phone_148,wall_21]=True
  close_item[phone_148,microwave_86]=True
  close_item[phone_148,wall_150]=True
  close_item[phone_148,light_187]=True
  close_item[phone_148,wall_28]=True
  inside[ceiling_326,home_office_248]=True
  close_item[napkin_2019,cupboard_64]=True
  inside[hanger_264,home_office_248]=True
  inside[hanger_264,dresser_258]=True
  close_item[kitchen_counter_1000,knife_2017]=True
  on[cupboard_65,wall_21]=True
  on[ceiling_154,wall_151]=True
  close_item[toilet_166,floor_160]=True
  close_item[toilet_166,floor_161]=True
  close_item[toilet_166,doorjamb_32]=True
  close_item[toilet_166,floor_2]=True
  close_item[toilet_166,floor_3]=True
  close_item[toilet_166,floor_6]=True
  close_item[toilet_166,shower_167]=True
  close_item[toilet_166,mat_135]=True
  close_item[toilet_166,shower_169]=True
  close_item[toilet_166,curtain_170]=True
  close_item[toilet_166,freezer_80]=True
  close_item[toilet_166,light_146]=True
  close_item[toilet_166,powersocket_147]=True
  close_item[toilet_166,wall_150]=True
  close_item[toilet_166,wall_22]=True
  close_item[toilet_166,wall_153]=True
  close_item[toilet_166,wall_28]=True
  close_item[toilet_166,door_31]=True
  close_item[bathroom_counter_171,floor_162]=True
  close_item[bathroom_counter_171,walllamp_163]=True
  close_item[bathroom_counter_171,walllamp_165]=True
  close_item[bathroom_counter_171,band_aids_2055]=True
  close_item[bathroom_counter_171,bathroom_cabinet_168]=True
  close_item[bathroom_counter_171,faucet_172]=True
  close_item[bathroom_counter_171,sink_173]=True
  close_item[bathroom_counter_171,toothbrush_holder_2061]=True
  close_item[bathroom_counter_171,wall_151]=True
  close_item[bathroom_counter_171,wall_152]=True
  close_item[bathroom_counter_171,mat_185]=True
  close_item[bathroom_counter_171,sponge_2040]=True
  close_item[bathroom_counter_171,floor_158]=True
  close_item[bathroom_counter_171,floor_159]=True
  on[hanger_2014,couch_257]=True
  inside[cutting_board_2025,dining_room_1]=True
  inside[cpuscreen_274,home_office_248]=True
  close_item[chair_191,desk_192]=True
  close_item[chair_191,mat_230]=True
  close_item[chair_191,floor_234]=True
  close_item[chair_191,floor_235]=True
  close_item[chair_191,photoframe_204]=True
  close_item[chair_191,floor_236]=True
  close_item[chair_191,wall_243]=True
  close_item[chair_191,wall_244]=True
  close_item[chair_191,wall_245]=True
  close_item[chair_191,wall_246]=True
  close_item[chair_191,bookshelf_190]=True
  close_item[light_196,wall_320]=True
  close_item[light_196,filing_cabinet_195]=True
  close_item[light_196,wall_323]=True
  close_item[light_196,mat_281]=True
  close_item[light_196,ceiling_327]=True
  close_item[light_196,ceiling_326]=True
  close_item[light_196,floor_237]=True
  close_item[light_196,floor_335]=True
  close_item[light_196,floor_336]=True
  close_item[light_196,ceiling_241]=True
  close_item[light_196,floor_337]=True
  close_item[light_196,wall_246]=True
  close_item[light_196,powersocket_279]=True
  close_item[light_196,light_280]=True
  close_item[light_196,doorjamb_345]=True
  close_item[light_196,door_347]=True
  close_item[light_196,bookshelf_253]=True
  inside[wallshelf_74,dining_room_1]=True
  inside[needle_2009,filing_cabinet_195]=True
  inside[needle_2009,bedroom_189]=True
  inside[floor_335,home_office_248]=True
  facing_item[ceiling_155,drawing_186]=True
  facing_item[chair_254,computer_273]=True
  inside[ceiling_242,bedroom_189]=True
  inside[drawing_283,home_office_248]=True
  facing_item[wall_22,drawing_139]=True
  facing_item[wall_22,drawing_140]=True
  facing_item[wall_22,drawing_141]=True
  facing_item[wall_22,drawing_142]=True
  on[ceiling_328,wall_322]=True
  inside[wall_319,home_office_248]=True
  on[kitchen_counter_70,floor_10]=True
  close_item[floor_161,floor_160]=True
  close_item[floor_161,floor_162]=True
  close_item[floor_161,mat_185]=True
  close_item[floor_161,photoframe_133]=True
  close_item[floor_161,toilet_166]=True
  close_item[floor_161,shower_167]=True
  close_item[floor_161,floor_6]=True
  close_item[floor_161,shower_169]=True
  close_item[floor_161,curtain_170]=True
  close_item[floor_161,nightstand_73]=True
  close_item[floor_161,freezer_80]=True
  close_item[floor_161,light_146]=True
  close_item[floor_161,powersocket_147]=True
  close_item[floor_161,wall_150]=True
  close_item[floor_161,wall_22]=True
  close_item[floor_161,wall_152]=True
  close_item[floor_161,wall_153]=True
  close_item[floor_161,door_31]=True
  facing_item[light_280,computer_273]=True
  facing_item[light_280,drawing_283]=True
  inside[tray_83,dining_room_1]=True
  inside[tray_83,oven_82]=True
  on[food_food_2045,plate_1004]=True
  close_item[drawing_186,floor_162]=True
  close_item[drawing_186,walllamp_165]=True
  close_item[drawing_186,wall_152]=True
  close_item[drawing_186,wall_153]=True
  close_item[drawing_186,ceiling_156]=True
  close_item[drawing_186,ceiling_157]=True
  inside[food_carrot_2018,bedroom_189]=True
  inside[closetdrawer_267,home_office_248]=True
  inside[closetdrawer_267,dresser_258]=True
  close_item[mat_230,desk_192]=True
  close_item[mat_230,nightstand_193]=True
  close_item[mat_230,bed_194]=True
  close_item[mat_230,door_229]=True
  close_item[mat_230,powersocket_197]=True
  close_item[mat_230,pillow_231]=True
  close_item[mat_230,floor_234]=True
  close_item[mat_230,floor_235]=True
  close_item[mat_230,floor_236]=True
  close_item[mat_230,photoframe_204]=True
  close_item[mat_230,floor_238]=True
  close_item[mat_230,floor_237]=True
  close_item[mat_230,toy_2034]=True
  close_item[mat_230,wall_243]=True
  close_item[mat_230,wall_244]=True
  close_item[mat_230,wall_245]=True
  close_item[mat_230,wall_246]=True
  close_item[mat_230,shoe_rack_2013]=True
  close_item[mat_230,bookshelf_190]=True
  close_item[mat_230,chair_191]=True
  inside[clothes_hat_2028,dining_room_1]=True
  facing_item[curtain_286,television_278]=True
  close_item[floor_234,nightstand_193]=True
  close_item[floor_234,bed_194]=True
  close_item[floor_234,doorjamb_228]=True
  close_item[floor_234,door_229]=True
  close_item[floor_234,powersocket_197]=True
  close_item[floor_234,mat_230]=True
  close_item[floor_234,pillow_231]=True
  close_item[floor_234,nightstand_72]=True
  close_item[floor_234,orchid_136]=True
  close_item[floor_234,floor_235]=True
  close_item[floor_234,photoframe_204]=True
  close_item[floor_234,floor_236]=True
  close_item[floor_234,floor_238]=True
  close_item[floor_234,floor_8]=True
  close_item[floor_234,wall_243]=True
  close_item[floor_234,wall_244]=True
  close_item[floor_234,wall_245]=True
  close_item[floor_234,wall_30]=True
  close_item[floor_234,bookshelf_190]=True
  close_item[floor_234,chair_191]=True
  on[ceiling_155,wall_150]=True
  inside[floor_338,home_office_248]=True
  inside[desk_251,home_office_248]=True
  close_item[nightstand_255,couch_256]=True
  close_item[nightstand_255,pillow_289]=True
  close_item[nightstand_255,pillow_288]=True
  close_item[nightstand_255,couch_257]=True
  close_item[nightstand_255,wall_324]=True
  close_item[nightstand_255,wall_323]=True
  close_item[nightstand_255,floor_335]=True
  close_item[nightstand_255,floor_336]=True
  close_item[nightstand_255,floor_341]=True
  close_item[nightstand_255,floor_342]=True
  close_item[nightstand_255,walllamp_314]=True
  close_item[nightstand_255,drawing_283]=True
  close_item[nightstand_255,tablelamp_317]=True
  close_item[nightstand_255,wall_318]=True
  facing_item[ceilinglamp_310,computer_273]=True
  facing_item[ceilinglamp_310,drawing_283]=True
  inside[walllamp_312,home_office_248]=True
  facing_item[ceilinglamp_164,drawing_186]=True
  close_item[oven_mitts_2005,filing_cabinet_195]=True
  inside[floor_5,dining_room_1]=True
  facing_item[floor_5,drawing_139]=True
  facing_item[floor_5,drawing_140]=True
  facing_item[floor_5,drawing_141]=True
  facing_item[floor_5,drawing_142]=True
  close_item[cup_2010,desk_251]=True
  inside[bookmark_2053,bedroom_189]=True
  close_item[food_food_2016,cupboard_65]=True
  inside[mousepad_276,home_office_248]=True
  on[toy_2034,mat_230]=True
  close_item[floor_162,floor_161]=True
  close_item[floor_162,wall_153]=True
  close_item[floor_162,walllamp_165]=True
  close_item[floor_162,bathroom_counter_171]=True
  close_item[floor_162,faucet_172]=True
  close_item[floor_162,sink_173]=True
  close_item[floor_162,wall_151]=True
  close_item[floor_162,wall_152]=True
  close_item[floor_162,mat_185]=True
  close_item[floor_162,drawing_186]=True
  close_item[floor_162,floor_158]=True
  close_item[floor_162,floor_159]=True
  on[clothes_shirt_2038,couch_256]=True
  close_item[hanger_261,wall_321]=True
  close_item[hanger_261,dresser_258]=True
  close_item[hanger_261,hanger_259]=True
  close_item[hanger_261,hanger_260]=True
  close_item[hanger_261,wall_325]=True
  close_item[hanger_261,hanger_262]=True
  close_item[hanger_261,hanger_263]=True
  close_item[hanger_261,hanger_264]=True
  close_item[hanger_261,hanger_265]=True
  close_item[hanger_261,closetdrawer_266]=True
  close_item[hanger_261,closetdrawer_267]=True
  close_item[hanger_261,closetdrawer_268]=True
  close_item[hanger_261,closetdrawer_269]=True
  close_item[hanger_261,ceiling_334]=True
  close_item[hanger_261,closetdrawer_270]=True
  close_item[hanger_261,ceiling_333]=True
  close_item[hanger_261,doorjamb_346]=True
  close_item[hanger_261,walllamp_315]=True
  inside[soap_2037,bathroom_149]=True
  inside[soap_2037,sink_173]=True
  inside[curtain_286,home_office_248]=True
  facing_item[floor_339,computer_273]=True
  close_item[walllamp_312,wall_325]=True
  close_item[walllamp_312,ceiling_329]=True
  close_item[walllamp_312,ceiling_334]=True
  close_item[walllamp_312,computer_273]=True
  close_item[walllamp_312,cpuscreen_274]=True
  close_item[walllamp_312,keyboard_275]=True
  close_item[walllamp_312,mousepad_276]=True
  close_item[walllamp_312,mouse_277]=True
  close_item[walllamp_312,floor_339]=True
  close_item[walllamp_312,desk_251]=True
  close_item[walllamp_312,wall_319]=True
  close_item[wall_245,light_280]=True
  close_item[wall_245,bookshelf_190]=True
  close_item[wall_245,chair_191]=True
  close_item[wall_245,desk_192]=True
  close_item[wall_245,wall_320]=True
  close_item[wall_245,wall_322]=True
  close_item[wall_245,filing_cabinet_195]=True
  close_item[wall_245,ceiling_328]=True
  close_item[wall_245,photoframe_204]=True
  close_item[wall_245,floor_338]=True
  close_item[wall_245,doorjamb_345]=True
  close_item[wall_245,door_347]=True
  close_item[wall_245,mat_230]=True
  close_item[wall_245,ceilinglamp_233]=True
  close_item[wall_245,floor_234]=True
  close_item[wall_245,floor_235]=True
  close_item[wall_245,floor_236]=True
  close_item[wall_245,floor_237]=True
  close_item[wall_245,ceiling_239]=True
  close_item[wall_245,ceiling_240]=True
  close_item[wall_245,ceiling_241]=True
  close_item[wall_245,wall_243]=True
  close_item[wall_245,wall_246]=True
  close_item[wall_245,bookshelf_250]=True
  inside[ceiling_14,dining_room_1]=True
  inside[basket_for_clothes_2062,home_office_248]=True
  inside[ceilinglamp_34,dining_room_1]=True
  facing_item[tablelamp_317,drawing_283]=True
  facing_item[tablelamp_317,television_278]=True
  close_item[ceiling_17,ceilinglamp_34]=True
  close_item[ceiling_17,shower_167]=True
  close_item[ceiling_17,shower_169]=True
  close_item[ceiling_17,drawing_139]=True
  close_item[ceiling_17,drawing_140]=True
  close_item[ceiling_17,drawing_141]=True
  close_item[ceiling_17,drawing_142]=True
  close_item[ceiling_17,ceiling_14]=True
  close_item[ceiling_17,freezer_80]=True
  close_item[ceiling_17,ceiling_16]=True
  close_item[ceiling_17,light_146]=True
  close_item[ceiling_17,wall_22]=True
  close_item[ceiling_17,wall_153]=True
  close_item[ceiling_17,ceiling_156]=True
  close_item[food_food_2065,cupboard_64]=True
  facing_item[ceiling_329,computer_273]=True
  inside[chair_254,home_office_248]=True
  close_item[sponge_2029,kitchen_counter_69]=True
  close_item[hanger_263,dresser_258]=True
  close_item[hanger_263,hanger_259]=True
  close_item[hanger_263,hanger_260]=True
  close_item[hanger_263,hanger_261]=True
  close_item[hanger_263,hanger_262]=True
  close_item[hanger_263,wall_325]=True
  close_item[hanger_263,hanger_264]=True
  close_item[hanger_263,hanger_265]=True
  close_item[hanger_263,closetdrawer_266]=True
  close_item[hanger_263,closetdrawer_267]=True
  close_item[hanger_263,closetdrawer_268]=True
  close_item[hanger_263,closetdrawer_269]=True
  close_item[hanger_263,ceiling_334]=True
  close_item[hanger_263,closetdrawer_270]=True
  close_item[hanger_263,doorjamb_346]=True
  close_item[hanger_263,walllamp_315]=True
  inside[kitchen_counter_69,dining_room_1]=True
  close_item[closetdrawer_268,dresser_258]=True
  close_item[closetdrawer_268,hanger_259]=True
  close_item[closetdrawer_268,hanger_260]=True
  close_item[closetdrawer_268,hanger_261]=True
  close_item[closetdrawer_268,hanger_262]=True
  close_item[closetdrawer_268,hanger_263]=True
  close_item[closetdrawer_268,closetdrawer_266]=True
  close_item[closetdrawer_268,closetdrawer_267]=True
  close_item[closetdrawer_268,closetdrawer_269]=True
  close_item[closetdrawer_268,closetdrawer_270]=True
  close_item[closetdrawer_268,closetdrawer_271]=True
  close_item[closetdrawer_268,closetdrawer_272]=True
  close_item[closetdrawer_268,television_278]=True
  close_item[closetdrawer_268,curtain_284]=True
  close_item[closetdrawer_268,curtain_285]=True
  close_item[closetdrawer_268,walllamp_315]=True
  close_item[closetdrawer_268,wall_321]=True
  close_item[closetdrawer_268,wall_325]=True
  close_item[closetdrawer_268,floor_343]=True
  close_item[closetdrawer_268,floor_344]=True
  close_item[closetdrawer_268,window_348]=True
  close_item[closetdrawer_268,tvstand_252]=True
  inside[dish_soap_1006,dishwasher_1002]=True
  inside[dish_soap_1006,bedroom_189]=True
  facing_item[wallshelf_74,drawing_138]=True
  facing_item[wallshelf_74,drawing_139]=True
  facing_item[wallshelf_74,drawing_140]=True
  facing_item[wallshelf_74,drawing_141]=True
  inside[toilet_166,bathroom_149]=True
  inside[toilet_166,shower_167]=True
  inside[kitchen_counter_1000,bedroom_189]=True
  inside[ceiling_17,dining_room_1]=True
  inside[food_food_2065,cupboard_64]=True
  inside[food_food_2065,dining_room_1]=True
  on[bookshelf_250,floor_338]=True
  close_item[tvstand_252,wall_321]=True
  close_item[tvstand_252,dresser_258]=True
  close_item[tvstand_252,wall_325]=True
  close_item[tvstand_252,closetdrawer_267]=True
  close_item[tvstand_252,closetdrawer_268]=True
  close_item[tvstand_252,closetdrawer_271]=True
  close_item[tvstand_252,floor_339]=True
  close_item[tvstand_252,window_348]=True
  close_item[tvstand_252,floor_340]=True
  close_item[tvstand_252,television_278]=True
  close_item[tvstand_252,floor_343]=True
  close_item[tvstand_252,floor_344]=True
  close_item[tvstand_252,table_249]=True
  close_item[tvstand_252,orchid_282]=True
  close_item[tvstand_252,walllamp_315]=True
  close_item[tvstand_252,curtain_284]=True
  close_item[tvstand_252,curtain_285]=True
  inside[floor_237,bedroom_189]=True
  facing_item[wall_152,drawing_186]=True
  inside[clothes_underwear_2049,home_office_248]=True
  close_item[floor_158,floor_160]=True
  close_item[floor_158,floor_162]=True
  close_item[floor_158,walllamp_163]=True
  close_item[floor_158,bathroom_counter_171]=True
  close_item[floor_158,faucet_172]=True
  close_item[floor_158,sink_173]=True
  close_item[floor_158,wall_150]=True
  close_item[floor_158,wall_151]=True
  close_item[floor_158,wall_152]=True
  close_item[floor_158,mat_185]=True
  close_item[floor_158,floor_159]=True
  inside[hanger_262,home_office_248]=True
  inside[hanger_262,dresser_258]=True
  close_item[walllamp_163,bathroom_cabinet_168]=True
  close_item[walllamp_163,bathroom_counter_171]=True
  close_item[walllamp_163,wall_151]=True
  close_item[walllamp_163,ceiling_154]=True
  close_item[walllamp_163,floor_158]=True
  close_item[walllamp_163,floor_159]=True
  close_item[dresser_258,hanger_259]=True
  close_item[dresser_258,hanger_260]=True
  close_item[dresser_258,hanger_261]=True
  close_item[dresser_258,hanger_262]=True
  close_item[dresser_258,hanger_263]=True
  close_item[dresser_258,hanger_264]=True
  close_item[dresser_258,hanger_265]=True
  close_item[dresser_258,closetdrawer_266]=True
  close_item[dresser_258,closetdrawer_267]=True
  close_item[dresser_258,closetdrawer_268]=True
  close_item[dresser_258,closetdrawer_269]=True
  close_item[dresser_258,closetdrawer_270]=True
  close_item[dresser_258,closetdrawer_271]=True
  close_item[dresser_258,closetdrawer_272]=True
  close_item[dresser_258,basket_for_clothes_2058]=True
  close_item[dresser_258,shoes_2066]=True
  close_item[dresser_258,television_278]=True
  close_item[dresser_258,curtain_284]=True
  close_item[dresser_258,curtain_285]=True
  close_item[dresser_258,walllamp_315]=True
  close_item[dresser_258,wall_321]=True
  close_item[dresser_258,wall_325]=True
  close_item[dresser_258,ceiling_334]=True
  close_item[dresser_258,floor_344]=True
  close_item[dresser_258,doorjamb_346]=True
  close_item[dresser_258,window_348]=True
  close_item[dresser_258,sheets_2043]=True
  close_item[dresser_258,tvstand_252]=True
  on[cup_2010,desk_251]=True
  inside[shower_169,bathroom_149]=True
  on[bathroom_cabinet_168,wall_151]=True
  inside[floor_10,dining_room_1]=True
  facing_item[mat_281,computer_273]=True
  facing_item[mat_281,drawing_283]=True
  close_item[ceiling_327,wall_320]=True
  close_item[ceiling_327,wall_322]=True
  close_item[ceiling_327,wall_323]=True
  close_item[ceiling_327,light_196]=True
  close_item[ceiling_327,ceiling_326]=True
  close_item[ceiling_327,ceiling_328]=True
  close_item[ceiling_327,ceiling_330]=True
  close_item[ceiling_327,ceiling_241]=True
  close_item[ceiling_327,ceilinglamp_310]=True
  close_item[ceiling_327,wall_246]=True
  close_item[ceiling_327,light_280]=True
  close_item[ceiling_327,doorjamb_345]=True
  close_item[ceiling_327,bookshelf_250]=True
  close_item[ceiling_327,bookshelf_253]=True
  inside[photoframe_133,dining_room_1]=True
  close_item[floor_342,pillow_288]=True
  close_item[floor_342,couch_257]=True
  close_item[floor_342,pillow_290]=True
  close_item[floor_342,pillow_289]=True
  close_item[floor_342,wall_324]=True
  close_item[floor_342,couch_256]=True
  close_item[floor_342,pillow_287]=True
  close_item[floor_342,floor_341]=True
  close_item[floor_342,floor_343]=True
  close_item[floor_342,table_249]=True
  close_item[floor_342,orchid_282]=True
  close_item[floor_342,walllamp_316]=True
  close_item[floor_342,tablelamp_317]=True
  close_item[floor_342,nightstand_255]=True
  inside[basket_for_clothes_2058,home_office_248]=True
  inside[basket_for_clothes_2058,dresser_258]=True
  inside[mat_230,bedroom_189]=True
  close_item[chair_60,ceilinglamp_35]=True
  close_item[chair_60,floor_4]=True
  close_item[chair_60,floor_5]=True
  close_item[chair_60,floor_7]=True
  close_item[chair_60,floor_8]=True
  close_item[chair_60,wall_30]=True
  close_item[chair_60,chair_59]=True
  close_item[chair_60,chair_61]=True
  close_item[chair_60,chair_62]=True
  close_item[chair_60,table_63]=True
  on[band_aids_2055,bathroom_counter_171]=True
  close_item[wall_153,photoframe_133]=True
  close_item[wall_153,floor_6]=True
  close_item[wall_153,ceiling_17]=True
  close_item[wall_153,light_146]=True
  close_item[wall_153,powersocket_147]=True
  close_item[wall_153,wall_150]=True
  close_item[wall_153,wall_22]=True
  close_item[wall_153,wall_152]=True
  close_item[wall_153,ceiling_155]=True
  close_item[wall_153,wall_28]=True
  close_item[wall_153,ceiling_156]=True
  close_item[wall_153,ceiling_157]=True
  close_item[wall_153,door_31]=True
  close_item[wall_153,floor_160]=True
  close_item[wall_153,floor_161]=True
  close_item[wall_153,floor_162]=True
  close_item[wall_153,doorjamb_32]=True
  close_item[wall_153,ceilinglamp_164]=True
  close_item[wall_153,toilet_166]=True
  close_item[wall_153,shower_167]=True
  close_item[wall_153,shower_169]=True
  close_item[wall_153,curtain_170]=True
  close_item[wall_153,mat_185]=True
  close_item[wall_153,drawing_186]=True
  close_item[wall_153,nightstand_73]=True
  close_item[wall_153,freezer_80]=True
  on[desk_251,floor_339]=True
  on[cup_1001,kitchen_counter_1000]=True
  inside[drawing_142,dining_room_1]=True
  facing_item[walllamp_165,drawing_186]=True
  inside[floor_162,bathroom_149]=True
  inside[ceilinglamp_233,bedroom_189]=True
  close_item[food_food_2008,table_249]=True
  inside[ceiling_330,home_office_248]=True
  facing_item[closetdrawer_267,computer_273]=True
  inside[powersocket_197,bedroom_189]=True
  on[ceiling_240,wall_245]=True
  close_item[ceiling_154,walllamp_163]=True
  close_item[ceiling_154,ceilinglamp_164]=True
  close_item[ceiling_154,bathroom_cabinet_168]=True
  close_item[ceiling_154,faucet_172]=True
  close_item[ceiling_154,wall_150]=True
  close_item[ceiling_154,wall_151]=True
  close_item[ceiling_154,wall_152]=True
  close_item[ceiling_154,ceiling_155]=True
  close_item[ceiling_154,ceiling_157]=True
  close_item[floor_160,doorjamb_32]=True
  close_item[floor_160,floor_161]=True
  close_item[floor_160,floor_159]=True
  close_item[floor_160,floor_2]=True
  close_item[floor_160,floor_3]=True
  close_item[floor_160,wall_153]=True
  close_item[floor_160,toilet_166]=True
  close_item[floor_160,shower_167]=True
  close_item[floor_160,mat_135]=True
  close_item[floor_160,freezer_80]=True
  close_item[floor_160,light_146]=True
  close_item[floor_160,powersocket_147]=True
  close_item[floor_160,wall_150]=True
  close_item[floor_160,wall_151]=True
  close_item[floor_160,mat_185]=True
  close_item[floor_160,light_187]=True
  close_item[floor_160,wall_28]=True
  close_item[floor_160,floor_158]=True
  close_item[floor_160,door_31]=True
  close_item[pot_98,cupboard_64]=True
  close_item[pot_98,pot_97]=True
  close_item[pot_98,kitchen_counter_66]=True
  close_item[pot_98,cupboard_65]=True
  close_item[pot_98,walllamp_36]=True
  close_item[pot_98,kitchen_counter_69]=True
  close_item[pot_98,floor_11]=True
  close_item[pot_98,toaster_76]=True
  close_item[pot_98,ceiling_12]=True
  close_item[pot_98,stovefan_79]=True
  close_item[pot_98,dishwasher_81]=True
  close_item[pot_98,oven_82]=True
  close_item[pot_98,tray_83]=True
  close_item[pot_98,wall_21]=True
  close_item[pot_98,wall_24]=True
  close_item[pot_98,wall_25]=True
  close_item[pot_98,wall_26]=True
  close_item[pot_98,knifeblock_92]=True
  close_item[pot_98,wall_29]=True
  inside[curtain_145,dining_room_1]=True
  on[desk_192,floor_236]=True
  on[ceiling_326,wall_323]=True
  on[ceiling_156,wall_153]=True
  inside[floor_339,home_office_248]=True
  on[dog_2000,couch_71]=True
  close_item[floor_9,kitchen_counter_66]=True
  close_item[floor_9,sink_67]=True
  close_item[floor_9,faucet_68]=True
  close_item[floor_9,floor_2]=True
  close_item[floor_9,floor_3]=True
  close_item[floor_9,mat_135]=True
  close_item[floor_9,floor_11]=True
  close_item[floor_9,toaster_76]=True
  close_item[floor_9,oven_82]=True
  close_item[floor_9,tray_83]=True
  close_item[floor_9,phone_148]=True
  close_item[floor_9,wall_21]=True
  close_item[floor_9,microwave_86]=True
  close_item[floor_9,wall_24]=True
  close_item[floor_9,light_187]=True
  close_item[floor_9,chair_61]=True
  close_item[floor_9,door_31]=True
  close_item[keyboard_2057,desk_251]=True
  on[cpuscreen_274,desk_251]=True
  on[door_31,floor_2]=True
  on[door_31,floor_3]=True
  close_item[clothes_scarf_2004,couch_71]=True
  on[television_278,tvstand_252]=True
  on[ceiling_19,wall_29]=True
  facing_item[floor_2,drawing_139]=True
  facing_item[floor_2,drawing_140]=True
  facing_item[floor_2,drawing_141]=True
  facing_item[floor_2,drawing_142]=True
  facing_item[mousepad_276,computer_273]=True
  on[wooden_spoon_2067,kitchen_counter_70]=True
  inside[bookshelf_190,bedroom_189]=True
  close_item[sink_173,floor_162]=True
  close_item[sink_173,bathroom_cabinet_168]=True
  close_item[sink_173,bathroom_counter_171]=True
  close_item[sink_173,faucet_172]=True
  close_item[sink_173,soap_2037]=True
  close_item[sink_173,wall_151]=True
  close_item[sink_173,wall_152]=True
  close_item[sink_173,mat_185]=True
  close_item[sink_173,floor_158]=True
  close_item[sink_173,floor_159]=True
  on[ceiling_239,wall_243]=True
  close_item[hanger_260,dresser_258]=True
  close_item[hanger_260,hanger_259]=True
  close_item[hanger_260,hanger_261]=True
  close_item[hanger_260,hanger_262]=True
  close_item[hanger_260,hanger_263]=True
  close_item[hanger_260,hanger_264]=True
  close_item[hanger_260,hanger_265]=True
  close_item[hanger_260,closetdrawer_266]=True
  close_item[hanger_260,closetdrawer_267]=True
  close_item[hanger_260,closetdrawer_268]=True
  close_item[hanger_260,closetdrawer_269]=True
  close_item[hanger_260,closetdrawer_270]=True
  close_item[hanger_260,curtain_284]=True
  close_item[hanger_260,curtain_285]=True
  close_item[hanger_260,walllamp_315]=True
  close_item[hanger_260,wall_321]=True
  close_item[hanger_260,wall_325]=True
  close_item[hanger_260,ceiling_333]=True
  close_item[hanger_260,ceiling_334]=True
  close_item[hanger_260,doorjamb_346]=True
  close_item[hanger_260,window_348]=True
  close_item[keyboard_275,wall_322]=True
  close_item[keyboard_275,computer_273]=True
  close_item[keyboard_275,cpuscreen_274]=True
  close_item[keyboard_275,floor_339]=True
  close_item[keyboard_275,mousepad_276]=True
  close_item[keyboard_275,mouse_277]=True
  close_item[keyboard_275,floor_338]=True
  close_item[keyboard_275,walllamp_311]=True
  close_item[keyboard_275,walllamp_312]=True
  close_item[keyboard_275,desk_251]=True
  close_item[keyboard_275,chair_254]=True
  close_item[keyboard_275,wall_319]=True
  inside[pot_97,dining_room_1]=True
  inside[drawing_138,dining_room_1]=True
  facing_item[wall_153,drawing_186]=True
  facing_item[floor_336,drawing_283]=True
  inside[sheets_2032,bedroom_189]=True
  inside[chair_61,dining_room_1]=True
  close_item[wall_244,nightstand_193]=True
  close_item[wall_244,bed_194]=True
  close_item[wall_244,doorjamb_228]=True
  close_item[wall_244,door_229]=True
  close_item[wall_244,mat_230]=True
  close_item[wall_244,pillow_231]=True
  close_item[wall_244,pillow_232]=True
  close_item[wall_244,ceilinglamp_233]=True
  close_item[wall_244,floor_234]=True
  close_item[wall_244,floor_235]=True
  close_item[wall_244,floor_237]=True
  close_item[wall_244,floor_238]=True
  close_item[wall_244,ceiling_239]=True
  close_item[wall_244,ceiling_241]=True
  close_item[wall_244,ceiling_242]=True
  close_item[wall_244,wall_243]=True
  close_item[wall_244,wall_246]=True
  close_item[wall_244,chair_191]=True
  on[dvd_player_2047,table_249]=True
  close_item[floor_11,pot_97]=True
  close_item[floor_11,pot_98]=True
  close_item[floor_11,kitchen_counter_66]=True
  close_item[floor_11,sink_67]=True
  close_item[floor_11,kitchen_counter_69]=True
  close_item[floor_11,floor_4]=True
  close_item[floor_11,faucet_68]=True
  close_item[floor_11,floor_9]=True
  close_item[floor_11,floor_10]=True
  close_item[floor_11,toaster_76]=True
  close_item[floor_11,dishwasher_81]=True
  close_item[floor_11,oven_82]=True
  close_item[floor_11,tray_83]=True
  close_item[floor_11,wall_29]=True
  close_item[floor_11,wall_21]=True
  close_item[floor_11,wall_26]=True
  close_item[floor_11,chair_61]=True
  close_item[floor_11,chair_62]=True
  close_item[floor_11,table_63]=True
  close_item[toothbrush_holder_2059,filing_cabinet_195]=True
  close_item[ceiling_16,ceilinglamp_34]=True
  close_item[ceiling_16,ceilinglamp_35]=True
  close_item[ceiling_16,couch_71]=True
  close_item[ceiling_16,drawing_138]=True
  close_item[ceiling_16,drawing_139]=True
  close_item[ceiling_16,drawing_140]=True
  close_item[ceiling_16,drawing_141]=True
  close_item[ceiling_16,drawing_142]=True
  close_item[ceiling_16,ceiling_15]=True
  close_item[ceiling_16,ceiling_17]=True
  close_item[ceiling_16,ceiling_20]=True
  close_item[ceiling_16,wall_22]=True
  close_item[ceiling_16,wall_23]=True
  close_item[ceiling_16,wall_30]=True
  close_item[walllamp_36,cupboard_64]=True
  close_item[walllamp_36,pot_97]=True
  close_item[walllamp_36,pot_98]=True
  close_item[walllamp_36,cupboard_65]=True
  close_item[walllamp_36,kitchen_counter_66]=True
  close_item[walllamp_36,kitchen_counter_69]=True
  close_item[walllamp_36,toaster_76]=True
  close_item[walllamp_36,ceiling_12]=True
  close_item[walllamp_36,ceiling_13]=True
  close_item[walllamp_36,stovefan_79]=True
  close_item[walllamp_36,oven_82]=True
  close_item[walllamp_36,tray_83]=True
  close_item[walllamp_36,wall_21]=True
  close_item[walllamp_36,wall_24]=True
  close_item[walllamp_36,wall_25]=True
  close_item[walllamp_36,wall_26]=True
  close_item[walllamp_36,knifeblock_92]=True
  close_item[walllamp_36,wall_29]=True
  inside[floor_342,home_office_248]=True
  surfaces[floor_2] = True
  surfaces[floor_3] = True
  surfaces[floor_4] = True
  surfaces[floor_5] = True
  surfaces[floor_6] = True
  surfaces[floor_7] = True
  surfaces[floor_8] = True
  surfaces[floor_9] = True
  surfaces[floor_10] = True
  surfaces[floor_11] = True
  can_open[door_31] = True
  movable[chair_59] = True
  surfaces[chair_59] = True
  grabbable[chair_59] = True
  sittable[chair_59] = True
  movable[chair_60] = True
  surfaces[chair_60] = True
  grabbable[chair_60] = True
  sittable[chair_60] = True
  movable[chair_61] = True
  surfaces[chair_61] = True
  grabbable[chair_61] = True
  sittable[chair_61] = True
  movable[chair_62] = True
  surfaces[chair_62] = True
  grabbable[chair_62] = True
  sittable[chair_62] = True
  movable[table_63] = True
  surfaces[table_63] = True
  can_open[cupboard_64] = True
  containers[cupboard_64] = True
  can_open[cupboard_65] = True
  containers[cupboard_65] = True
  surfaces[kitchen_counter_66] = True
  recipient[sink_67] = True
  containers[sink_67] = True
  has_switch[faucet_68] = True
  surfaces[kitchen_counter_69] = True
  surfaces[kitchen_counter_70] = True
  movable[couch_71] = True
  surfaces[couch_71] = True
  lieable[couch_71] = True
  sittable[couch_71] = True
  surfaces[nightstand_72] = True
  can_open[nightstand_72] = True
  containers[nightstand_72] = True
  surfaces[nightstand_73] = True
  can_open[nightstand_73] = True
  containers[nightstand_73] = True
  has_switch[toaster_76] = True
  movable[toaster_76] = True
  has_plug[toaster_76] = True
  has_switch[freezer_80] = True
  has_plug[freezer_80] = True
  can_open[freezer_80] = True
  containers[freezer_80] = True
  has_switch[dishwasher_81] = True
  can_open[dishwasher_81] = True
  containers[dishwasher_81] = True
  has_switch[oven_82] = True
  has_plug[oven_82] = True
  can_open[oven_82] = True
  containers[oven_82] = True
  movable[tray_83] = True
  surfaces[tray_83] = True
  grabbable[tray_83] = True
  containers[coffe_maker_84] = True
  can_open[coffe_maker_84] = True
  has_switch[coffe_maker_84] = True
  has_plug[coffe_maker_84] = True
  movable[coffe_maker_84] = True
  recipient[coffe_maker_84] = True
  has_switch[microwave_86] = True
  has_plug[microwave_86] = True
  can_open[microwave_86] = True
  containers[microwave_86] = True
  movable[pot_97] = True
  recipient[pot_97] = True
  can_open[pot_97] = True
  grabbable[pot_97] = True
  movable[pot_98] = True
  recipient[pot_98] = True
  can_open[pot_98] = True
  grabbable[pot_98] = True
  grabbable[mat_135] = True
  sittable[mat_135] = True
  lieable[mat_135] = True
  surfaces[mat_135] = True
  movable[mat_135] = True
  cuttable[drawing_138] = True
  grabbable[drawing_138] = True
  lookable[drawing_138] = True
  movable[drawing_138] = True
  has_paper[drawing_138] = True
  cuttable[drawing_139] = True
  grabbable[drawing_139] = True
  lookable[drawing_139] = True
  movable[drawing_139] = True
  has_paper[drawing_139] = True
  cuttable[drawing_140] = True
  grabbable[drawing_140] = True
  lookable[drawing_140] = True
  movable[drawing_140] = True
  has_paper[drawing_140] = True
  cuttable[drawing_141] = True
  grabbable[drawing_141] = True
  lookable[drawing_141] = True
  movable[drawing_141] = True
  has_paper[drawing_141] = True
  cuttable[drawing_142] = True
  grabbable[drawing_142] = True
  lookable[drawing_142] = True
  movable[drawing_142] = True
  has_paper[drawing_142] = True
  movable[curtain_143] = True
  can_open[curtain_143] = True
  cover_object[curtain_143] = True
  movable[curtain_144] = True
  can_open[curtain_144] = True
  cover_object[curtain_144] = True
  movable[curtain_145] = True
  can_open[curtain_145] = True
  cover_object[curtain_145] = True
  has_switch[light_146] = True
  has_plug[light_146] = True
  has_switch[phone_148] = True
  movable[phone_148] = True
  has_plug[phone_148] = True
  grabbable[phone_148] = True
  surfaces[floor_158] = True
  surfaces[floor_159] = True
  surfaces[floor_160] = True
  surfaces[floor_161] = True
  surfaces[floor_162] = True
  can_open[toilet_166] = True
  sittable[toilet_166] = True
  containers[toilet_166] = True
  surfaces[bathroom_cabinet_168] = True
  can_open[bathroom_cabinet_168] = True
  containers[bathroom_cabinet_168] = True
  movable[curtain_170] = True
  can_open[curtain_170] = True
  cover_object[curtain_170] = True
  surfaces[bathroom_counter_171] = True
  has_switch[faucet_172] = True
  recipient[sink_173] = True
  containers[sink_173] = True
  grabbable[mat_185] = True
  sittable[mat_185] = True
  lieable[mat_185] = True
  surfaces[mat_185] = True
  movable[mat_185] = True
  cuttable[drawing_186] = True
  grabbable[drawing_186] = True
  lookable[drawing_186] = True
  movable[drawing_186] = True
  has_paper[drawing_186] = True
  has_switch[light_187] = True
  has_plug[light_187] = True
  surfaces[bookshelf_190] = True
  can_open[bookshelf_190] = True
  containers[bookshelf_190] = True
  movable[chair_191] = True
  surfaces[chair_191] = True
  grabbable[chair_191] = True
  sittable[chair_191] = True
  movable[desk_192] = True
  surfaces[desk_192] = True
  surfaces[nightstand_193] = True
  can_open[nightstand_193] = True
  containers[nightstand_193] = True
  surfaces[bed_194] = True
  lieable[bed_194] = True
  sittable[bed_194] = True
  surfaces[filing_cabinet_195] = True
  can_open[filing_cabinet_195] = True
  containers[filing_cabinet_195] = True
  has_switch[light_196] = True
  has_plug[light_196] = True
  can_open[door_229] = True
  grabbable[mat_230] = True
  sittable[mat_230] = True
  lieable[mat_230] = True
  surfaces[mat_230] = True
  movable[mat_230] = True
  movable[pillow_231] = True
  grabbable[pillow_231] = True
  movable[pillow_232] = True
  grabbable[pillow_232] = True
  surfaces[floor_234] = True
  surfaces[floor_235] = True
  surfaces[floor_236] = True
  surfaces[floor_237] = True
  surfaces[floor_238] = True
  movable[table_249] = True
  surfaces[table_249] = True
  surfaces[bookshelf_250] = True
  can_open[bookshelf_250] = True
  containers[bookshelf_250] = True
  movable[desk_251] = True
  surfaces[desk_251] = True
  surfaces[tvstand_252] = True
  surfaces[bookshelf_253] = True
  can_open[bookshelf_253] = True
  containers[bookshelf_253] = True
  movable[chair_254] = True
  surfaces[chair_254] = True
  grabbable[chair_254] = True
  sittable[chair_254] = True
  surfaces[nightstand_255] = True
  can_open[nightstand_255] = True
  containers[nightstand_255] = True
  movable[couch_256] = True
  surfaces[couch_256] = True
  lieable[couch_256] = True
  sittable[couch_256] = True
  movable[couch_257] = True
  surfaces[couch_257] = True
  lieable[couch_257] = True
  sittable[couch_257] = True
  can_open[dresser_258] = True
  containers[dresser_258] = True
  movable[hanger_259] = True
  grabbable[hanger_259] = True
  hangable[hanger_259] = True
  movable[hanger_260] = True
  grabbable[hanger_260] = True
  hangable[hanger_260] = True
  movable[hanger_261] = True
  grabbable[hanger_261] = True
  hangable[hanger_261] = True
  movable[hanger_262] = True
  grabbable[hanger_262] = True
  hangable[hanger_262] = True
  movable[hanger_263] = True
  grabbable[hanger_263] = True
  hangable[hanger_263] = True
  movable[hanger_264] = True
  grabbable[hanger_264] = True
  hangable[hanger_264] = True
  movable[hanger_265] = True
  grabbable[hanger_265] = True
  hangable[hanger_265] = True
  has_switch[computer_273] = True
  lookable[computer_273] = True
  movable[keyboard_275] = True
  has_plug[keyboard_275] = True
  grabbable[keyboard_275] = True
  movable[mousepad_276] = True
  surfaces[mousepad_276] = True
  movable[mouse_277] = True
  has_plug[mouse_277] = True
  grabbable[mouse_277] = True
  has_switch[television_278] = True
  has_plug[television_278] = True
  lookable[television_278] = True
  has_switch[light_280] = True
  has_plug[light_280] = True
  grabbable[mat_281] = True
  sittable[mat_281] = True
  lieable[mat_281] = True
  surfaces[mat_281] = True
  movable[mat_281] = True
  cuttable[drawing_283] = True
  grabbable[drawing_283] = True
  lookable[drawing_283] = True
  movable[drawing_283] = True
  has_paper[drawing_283] = True
  movable[curtain_284] = True
  can_open[curtain_284] = True
  cover_object[curtain_284] = True
  movable[curtain_285] = True
  can_open[curtain_285] = True
  cover_object[curtain_285] = True
  movable[curtain_286] = True
  can_open[curtain_286] = True
  cover_object[curtain_286] = True
  movable[pillow_287] = True
  grabbable[pillow_287] = True
  movable[pillow_288] = True
  grabbable[pillow_288] = True
  movable[pillow_289] = True
  grabbable[pillow_289] = True
  movable[pillow_290] = True
  grabbable[pillow_290] = True
  has_switch[tablelamp_317] = True
  surfaces[floor_335] = True
  surfaces[floor_336] = True
  surfaces[floor_337] = True
  surfaces[floor_338] = True
  surfaces[floor_339] = True
  surfaces[floor_340] = True
  surfaces[floor_341] = True
  surfaces[floor_342] = True
  surfaces[floor_343] = True
  surfaces[floor_344] = True
  can_open[door_347] = True
  surfaces[kitchen_counter_1000] = True
  movable[cup_1001] = True
  recipient[cup_1001] = True
  pourable[cup_1001] = True
  grabbable[cup_1001] = True
  has_switch[dishwasher_1002] = True
  can_open[dishwasher_1002] = True
  containers[dishwasher_1002] = True
  movable[cup_1003] = True
  recipient[cup_1003] = True
  pourable[cup_1003] = True
  grabbable[cup_1003] = True
  movable[plate_1004] = True
  surfaces[plate_1004] = True
  recipient[plate_1004] = True
  grabbable[plate_1004] = True
  movable[plate_1005] = True
  surfaces[plate_1005] = True
  recipient[plate_1005] = True
  grabbable[plate_1005] = True
  movable[dish_soap_1006] = True
  pourable[dish_soap_1006] = True
  grabbable[dish_soap_1006] = True
  cream[dish_soap_1006] = True
  movable[dog_2000] = True
  grabbable[dog_2000] = True
  movable[clothes_hat_2001] = True
  clothes[clothes_hat_2001] = True
  grabbable[clothes_hat_2001] = True
  hangable[clothes_hat_2001] = True
  grabbable[check_2002] = True
  movable[check_2002] = True
  has_paper[check_2002] = True
  readable[check_2002] = True
  grabbable[check_2003] = True
  movable[check_2003] = True
  has_paper[check_2003] = True
  readable[check_2003] = True
  movable[clothes_scarf_2004] = True
  clothes[clothes_scarf_2004] = True
  grabbable[clothes_scarf_2004] = True
  hangable[clothes_scarf_2004] = True
  movable[oven_mitts_2005] = True
  clothes[oven_mitts_2005] = True
  grabbable[oven_mitts_2005] = True
  hangable[oven_mitts_2005] = True
  movable[detergent_2006] = True
  pourable[detergent_2006] = True
  grabbable[detergent_2006] = True
  movable[clothes_dress_2007] = True
  clothes[clothes_dress_2007] = True
  grabbable[clothes_dress_2007] = True
  hangable[clothes_dress_2007] = True
  movable[food_food_2008] = True
  eatable[food_food_2008] = True
  grabbable[food_food_2008] = True
  cuttable[food_food_2008] = True
  movable[needle_2009] = True
  grabbable[needle_2009] = True
  movable[cup_2010] = True
  recipient[cup_2010] = True
  pourable[cup_2010] = True
  grabbable[cup_2010] = True
  movable[cd_2011] = True
  grabbable[cd_2011] = True
  movable[thread_2012] = True
  grabbable[thread_2012] = True
  cuttable[thread_2012] = True
  movable[shoe_rack_2013] = True
  surfaces[shoe_rack_2013] = True
  grabbable[shoe_rack_2013] = True
  movable[hanger_2014] = True
  grabbable[hanger_2014] = True
  hangable[hanger_2014] = True
  grabbable[form_2015] = True
  movable[form_2015] = True
  has_paper[form_2015] = True
  movable[food_food_2016] = True
  eatable[food_food_2016] = True
  grabbable[food_food_2016] = True
  cuttable[food_food_2016] = True
  movable[knife_2017] = True
  grabbable[knife_2017] = True
  movable[food_carrot_2018] = True
  eatable[food_carrot_2018] = True
  grabbable[food_carrot_2018] = True
  cuttable[food_carrot_2018] = True
  grabbable[napkin_2019] = True
  movable[napkin_2019] = True
  cover_object[napkin_2019] = True
  has_paper[napkin_2019] = True
  movable[soap_2020] = True
  grabbable[soap_2020] = True
  cream[soap_2020] = True
  movable[tray_2021] = True
  surfaces[tray_2021] = True
  grabbable[tray_2021] = True
  movable[food_peanut_butter_2022] = True
  eatable[food_peanut_butter_2022] = True
  grabbable[food_peanut_butter_2022] = True
  cream[food_peanut_butter_2022] = True
  movable[food_carrot_2023] = True
  eatable[food_carrot_2023] = True
  grabbable[food_carrot_2023] = True
  cuttable[food_carrot_2023] = True
  movable[knife_2024] = True
  grabbable[knife_2024] = True
  movable[cutting_board_2025] = True
  surfaces[cutting_board_2025] = True
  grabbable[cutting_board_2025] = True
  grabbable[juice_2026] = True
  movable[juice_2026] = True
  pourable[juice_2026] = True
  drinkable[juice_2026] = True
  grabbable[homework_2027] = True
  movable[homework_2027] = True
  has_paper[homework_2027] = True
  readable[homework_2027] = True
  movable[clothes_hat_2028] = True
  clothes[clothes_hat_2028] = True
  grabbable[clothes_hat_2028] = True
  hangable[clothes_hat_2028] = True
  movable[sponge_2029] = True
  grabbable[sponge_2029] = True
  movable[soap_2030] = True
  grabbable[soap_2030] = True
  cream[soap_2030] = True
  movable[food_food_2031] = True
  eatable[food_food_2031] = True
  grabbable[food_food_2031] = True
  cuttable[food_food_2031] = True
  grabbable[sheets_2032] = True
  movable[sheets_2032] = True
  cover_object[sheets_2032] = True
  movable[food_food_2033] = True
  eatable[food_food_2033] = True
  grabbable[food_food_2033] = True
  cuttable[food_food_2033] = True
  movable[toy_2034] = True
  grabbable[toy_2034] = True
  movable[food_butter_2035] = True
  grabbable[food_butter_2035] = True
  cream[food_butter_2035] = True
  movable[pasta_2036] = True
  pourable[pasta_2036] = True
  grabbable[pasta_2036] = True
  movable[soap_2037] = True
  grabbable[soap_2037] = True
  cream[soap_2037] = True
  movable[clothes_shirt_2038] = True
  clothes[clothes_shirt_2038] = True
  grabbable[clothes_shirt_2038] = True
  hangable[clothes_shirt_2038] = True
  movable[pencil_2039] = True
  grabbable[pencil_2039] = True
  movable[sponge_2040] = True
  grabbable[sponge_2040] = True
  movable[detergent_2041] = True
  pourable[detergent_2041] = True
  grabbable[detergent_2041] = True
  movable[food_orange_2042] = True
  eatable[food_orange_2042] = True
  grabbable[food_orange_2042] = True
  cuttable[food_orange_2042] = True
  grabbable[sheets_2043] = True
  movable[sheets_2043] = True
  cover_object[sheets_2043] = True
  movable[tea_bag_2044] = True
  grabbable[tea_bag_2044] = True
  movable[food_food_2045] = True
  eatable[food_food_2045] = True
  grabbable[food_food_2045] = True
  cuttable[food_food_2045] = True
  grabbable[bookmark_2046] = True
  movable[bookmark_2046] = True
  has_paper[bookmark_2046] = True
  can_open[dvd_player_2047] = True
  grabbable[dvd_player_2047] = True
  has_switch[dvd_player_2047] = True
  surfaces[dvd_player_2047] = True
  movable[dvd_player_2047] = True
  has_plug[dvd_player_2047] = True
  grabbable[form_2048] = True
  movable[form_2048] = True
  has_paper[form_2048] = True
  movable[clothes_underwear_2049] = True
  clothes[clothes_underwear_2049] = True
  grabbable[clothes_underwear_2049] = True
  hangable[clothes_underwear_2049] = True
  grabbable[coffee_filter_2050] = True
  movable[coffee_filter_2050] = True
  has_paper[coffee_filter_2050] = True
  readable[newspaper_2051] = True
  can_open[newspaper_2051] = True
  grabbable[newspaper_2051] = True
  has_paper[newspaper_2051] = True
  movable[newspaper_2051] = True
  cover_object[newspaper_2051] = True
  movable[clothes_socks_2052] = True
  clothes[clothes_socks_2052] = True
  grabbable[clothes_socks_2052] = True
  hangable[clothes_socks_2052] = True
  grabbable[bookmark_2053] = True
  movable[bookmark_2053] = True
  has_paper[bookmark_2053] = True
  grabbable[check_2054] = True
  movable[check_2054] = True
  has_paper[check_2054] = True
  readable[check_2054] = True
  movable[band_aids_2055] = True
  grabbable[band_aids_2055] = True
  cuttable[band_aids_2055] = True
  movable[detergent_2056] = True
  pourable[detergent_2056] = True
  grabbable[detergent_2056] = True
  movable[keyboard_2057] = True
  has_plug[keyboard_2057] = True
  grabbable[keyboard_2057] = True
  movable[basket_for_clothes_2058] = True
  can_open[basket_for_clothes_2058] = True
  grabbable[basket_for_clothes_2058] = True
  containers[basket_for_clothes_2058] = True
  movable[toothbrush_holder_2059] = True
  grabbable[toothbrush_holder_2059] = True
  containers[toothbrush_holder_2059] = True
  movable[ground_coffee_2060] = True
  can_open[ground_coffee_2060] = True
  grabbable[ground_coffee_2060] = True
  movable[toothbrush_holder_2061] = True
  grabbable[toothbrush_holder_2061] = True
  containers[toothbrush_holder_2061] = True
  movable[basket_for_clothes_2062] = True
  can_open[basket_for_clothes_2062] = True
  grabbable[basket_for_clothes_2062] = True
  containers[basket_for_clothes_2062] = True
  cream[after_shave_2063] = True
  can_open[after_shave_2063] = True
  grabbable[after_shave_2063] = True
  pourable[after_shave_2063] = True
  movable[after_shave_2063] = True
  movable[knife_2064] = True
  grabbable[knife_2064] = True
  movable[food_food_2065] = True
  eatable[food_food_2065] = True
  grabbable[food_food_2065] = True
  cuttable[food_food_2065] = True
  movable[shoes_2066] = True
  clothes[shoes_2066] = True
  grabbable[shoes_2066] = True
  movable[wooden_spoon_2067] = True
  grabbable[wooden_spoon_2067] = True
