domain "virtualhome"

typedef item: object
typedef character: object
typedef ObjectList: item[]

# Features without return type annotations are assumed to be returning boolean values.

#state
feature is_on(x: item)
feature is_off(x: item)
feature plugged(x: item)
feature unplugged(x: item)
feature open(x: item)
feature closed(x: item)
feature dirty(x: item)
feature clean(x: item)
feature sitting(x: character)
feature lying(x: character)
feature cut(x:item)
feature sleeping(x: character)

#relationship
feature on(x: item, y: item)
feature inside(x: item, y: item)
feature between(door: item, room: item)
feature close(x: item, y: item)
feature facing(x: item, y: item)

feature close_char(x: character, y: item)
feature facing_char(x: character, y: item)
feature inside_char(x: character, y: item)
feature on_char(x: character, y: item)
feature on_body(x:item, y: character)
feature holds_rh(x: character, y: item)
feature holds_lh(x: character, y: item)

#Properties
feature surfaces(x: item)
feature grabbable(x: item)
feature sittable(x: item)
feature lieable(x: item)
feature hangable(x: item)
feature drinkable(x: item)
feature eatable(x: item)
feature recipient(x: item)
feature cuttable(x: item)
feature pourable(x: item)
feature can_open(x: item)
feature has_switch(x: item)
feature readable(x: item)
feature lookable(x: item)
feature containers(x: item)
feature clothes(x: item)
feature person(x: item)
feature body_part(x: item)
feature cover_object(x: item)
feature has_plug(x: item)
feature has_paper(x: item)
feature movable(x: item)
feature cream(x: item)


object_constant char:character

#category
feature is_room(x: item)
feature is_comb(x:item)
feature is_pillow(x:item)
feature is_teeth(x:item)
feature is_face_soap(x:item)
feature is_sheets(x:item)
feature is_mail(x:item)
feature is_remote_control(x:item)
feature is_instrument_violin(x:item)
feature is_shoe_rack(x:item)
feature is_lighter(x:item)
feature is_food_vegetable(x:item)
feature is_phone(x:item)
feature is_table_cloth(x:item)
feature is_pajamas(x:item)
feature is_clothes_socks(x:item)
feature is_form(x:item)
feature is_face(x:item)
feature is_wall_clock(x:item)
feature is_food_egg(x:item)
feature is_printing_paper(x:item)
feature is_paper_towel(x:item)
feature is_legs_both(x:item)
feature is_glue(x:item)
feature is_towel(x:item)
feature is_coffee_table(x:item)
feature is_food_sugar(x:item)
feature is_microphone(x:item)
feature is_foundation(x:item)
feature is_curtain(x:item)
feature is_mouse(x:item)
feature is_duster(x:item)
feature is_food_turkey(x:item)
feature is_bookshelf(x:item)
feature is_clothes_pants(x:item)
feature is_food_onion(x:item)
feature is_table(x:item)
feature is_scrabble(x:item)
feature is_wallshelf(x:item)
feature is_sink(x:item)
feature is_controller(x:item)
feature is_instrument_piano(x:item)
feature is_food_snack(x:item)
feature is_coin(x:item)
feature is_tape(x:item)
feature is_thread(x:item)
feature is_towel_rack(x:item)
feature is_electrical_outlet(x:item)
feature is_dog(x:item)
feature is_bathroom(x:item)
feature is_hair(x:item)
feature is_oil(x:item)
feature is_sponge(x:item)
feature is_cd_player(x:item)
feature is_measuring_cup(x:item)
feature is_food_apple(x:item)
feature is_knifeblock(x:item)
feature is_tablelamp(x:item)
feature is_basket_for_clothes(x:item)
feature is_drinking_glass(x:item)
feature is_beer(x:item)
feature is_novel(x:item)
feature is_light_bulb(x:item)
feature is_bathroom_cabinet(x:item)
feature is_bench(x:item)
feature is_dirt(x:item)
feature is_food_orange(x:item)
feature is_clothes_jacket(x:item)
feature is_electric_shaver(x:item)
feature is_envelope(x:item)
feature is_coffee_cup(x:item)
feature is_cleaning_solution(x:item)
feature is_tea_bag(x:item)
feature is_dough(x:item)
feature is_longboard(x:item)
feature is_napkin(x:item)
feature is_clothes_skirt(x:item)
feature is_walllamp(x:item)
feature is_chef_knife(x:item)
feature is_video_game_controller(x:item)
feature is_detergent(x:item)
feature is_hairdryer(x:item)
feature is_balanceball(x:item)
feature is_mirror(x:item)
feature is_bedroom(x:item)
feature is_mop(x:item)
feature is_iron(x:item)
feature is_shoes(x:item)
feature is_cards(x:item)
feature is_bag(x:item)
feature is_fly(x:item)
feature is_toilet(x:item)
feature is_rag(x:item)
feature is_clothes_shirt(x:item)
feature is_fork(x:item)
feature is_woman(x:item)
feature is_closetdrawer(x:item)
feature is_laser_pointer(x:item)
feature is_deck_of_cards(x:item)
feature is_food_noodles(x:item)
feature is_razor(x:item)
feature is_hands_both(x:item)
feature is_dishrack(x:item)
feature is_cup(x:item)
feature is_console(x:item)
feature is_food_cheese(x:item)
feature is_video_game_console(x:item)
feature is_bathroom_counter(x:item)
feature is_kitchen_counter(x:item)
feature is_oven(x:item)
feature is_filing_cabinet(x:item)
feature is_plate(x:item)
feature is_brush(x:item)
feature is_toaster(x:item)
feature is_tooth_paste(x:item)
feature is_shoe_shine_kit(x:item)
feature is_pasta(x:item)
feature is_toothbrush(x:item)
feature is_keys(x:item)
feature is_shelf(x:item)
feature is_box(x:item)
feature is_standingmirror(x:item)
feature is_scissors(x:item)
feature is_board_game(x:item)
feature is_mop_bucket(x:item)
feature is_love_seat(x:item)
feature is_bed(x:item)
feature is_cloth_napkin(x:item)
feature is_sauce_pan(x:item)
feature is_drying_rack(x:item)
feature is_ceilingfan(x:item)
feature is_window(x:item)
feature is_photoframe(x:item)
feature is_facial_cleanser(x:item)
feature is_cd(x:item)
feature is_ceiling(x:item)
feature is_dining_room(x:item)
feature is_alarm_clock(x:item)
feature is_floor_lamp(x:item)
feature is_blender(x:item)
feature is_stovefan(x:item)
feature is_maindoor(x:item)
feature is_band_aids(x:item)
feature is_broom(x:item)
feature is_food_dessert(x:item)
feature is_food_bacon(x:item)
feature is_check(x:item)
feature is_diary(x:item)
feature is_kettle(x:item)
feature is_food_cake(x:item)
feature is_ceilinglamp(x:item)
feature is_bowl(x:item)
feature is_spoon(x:item)
feature is_chair(x:item)
feature is_clothes_dress(x:item)
feature is_dry_pasta(x:item)
feature is_pantry(x:item)
feature is_button(x:item)
feature is_needle(x:item)
feature is_food_donut(x:item)
feature is_coffee_filter(x:item)
feature is_piano_bench(x:item)
feature is_microwave(x:item)
feature is_food_bread(x:item)
feature is_door(x:item)
feature is_newspaper(x:item)
feature is_food_salt(x:item)
feature is_toilet_paper(x:item)
feature is_coffee_pot(x:item)
feature is_ground_coffee(x:item)
feature is_food_pizza(x:item)
feature is_headset(x:item)
feature is_food_peanut_butter(x:item)
feature is_man(x:item)
feature is_food_ice_cream(x:item)
feature is_laundry_detergent(x:item)
feature is_cpuscreen(x:item)
feature is_homework(x:item)
feature is_bookmark(x:item)
feature is_clothes_gloves(x:item)
feature is_toothbrush_holder(x:item)
feature is_ice(x:item)
feature is_doorjamb(x:item)
feature is_nightstand(x:item)
feature is_alcohol(x:item)
feature is_kitchen_cabinet(x:item)
feature is_food_fish(x:item)
feature is_food_steak(x:item)
feature is_dustpan(x:item)
feature is_colander(x:item)
feature is_washing_machine(x:item)
feature is_food_jam(x:item)
feature is_address_book(x:item)
feature is_tvstand(x:item)
feature is_dresser(x:item)
feature is_candle(x:item)
feature is_hanger(x:item)
feature is_milk(x:item)
feature is_food_carrot(x:item)
feature is_cupboard(x:item)
feature is_bathtub(x:item)
feature is_purse(x:item)
feature is_fax_machine(x:item)
feature is_cleaning_bottle(x:item)
feature is_tray(x:item)
feature is_garbage_can(x:item)
feature is_coffe_maker(x:item)
feature is_instrument_guitar(x:item)
feature is_food_food(x:item)
feature is_floor(x:item)
feature is_stamp(x:item)
feature is_crayon(x:item)
feature is_mousepad(x:item)
feature is_oven_mitts(x:item)
feature is_home_office(x:item)
feature is_jelly(x:item)
feature is_food_chicken(x:item)
feature is_nail_polish(x:item)
feature is_trashcan(x:item)
feature is_clothes_scarf(x:item)
feature is_cat(x:item)
feature is_ironing_board(x:item)
feature is_powersocket(x:item)
feature is_television(x:item)
feature is_desk(x:item)
feature is_food_cereal(x:item)
feature is_spectacles(x:item)
feature is_wine_glass(x:item)
feature is_faucet(x:item)
feature is_vacuum_cleaner(x:item)
feature is_chessboard(x:item)
feature is_child(x:item)
feature is_food_oatmeal(x:item)
feature is_dish_soap(x:item)
feature is_wooden_spoon(x:item)
feature is_shampoo(x:item)
feature is_dvd_player(x:item)
feature is_music_stand(x:item)
feature is_creditcard(x:item)
feature is_centerpiece(x:item)
feature is_food_rice(x:item)
feature is_wine(x:item)
feature is_couch(x:item)
feature is_computer(x:item)
feature is_orchid(x:item)
feature is_stereo(x:item)
feature is_vase(x:item)
feature is_shredder(x:item)
feature is_food_butter(x:item)
feature is_mouthwash(x:item)
feature is_after_shave(x:item)
feature is_clothes_underwear(x:item)
feature is_toy(x:item)
feature is_knife(x:item)
feature is_pot(x:item)
feature is_keyboard(x:item)
feature is_freezer(x:item)
feature is_coffee(x:item)
feature is_water_glass(x:item)
feature is_drawing(x:item)
feature is_shaving_cream(x:item)
feature is_blow_dryer(x:item)
feature is_soap(x:item)
feature is_shower(x:item)
feature is_picture(x:item)
feature is_clothes_hat(x:item)
feature is_wall(x:item)
feature is_cutting_board(x:item)
feature is_laptop(x:item)
feature is_arms_both(x:item)
feature is_pencil(x:item)
feature is_dishwasher(x:item)
feature is_food_kiwi(x:item)
feature is_water(x:item)
feature is_conditioner(x:item)
feature is_tea(x:item)
feature is_hairbrush(x:item)
feature is_feet_both(x:item)
feature is_mat(x:item)
feature is_juice(x:item)
feature is_light(x:item)
feature is_folder(x:item)
feature is_bills(x:item)


#controllers
controller walk_executor(x: item)
controller switchoff_executor(x: item)
controller switchon_executor(x: item)
controller put_executor(x: item, y: item)
controller grab_executor(x: item)
controller standup_executor(x: character)
controller wash_executor(x: item)
controller sit_executor(x: item)
controller lie_executor(x: item)
controller open_executor(x: item)
controller close_executor(x: item)
controller pour_executor(x: item, y: item)
controller plugin_executor(x: item)
controller plugout_executor(x: item)
controller find_executor(x: item)
controller turnto_executor(x: item)
controller cut_executor(x: item)
controller eat_executor(x: item)
controller sleep_executor(x: character)
controller greet_executor(x: item)
controller drink_executor(x: item)
controller lookat_executor(x: item)
controller wipe_executor(x: item)
controller puton_executor(x: item)
controller putoff_executor(x: item)
controller read_executor(x: item)
controller touch_executor(x: item)
controller type_executor(x: item)
controller watch_executor(x: item)
controller move_executor(x: item)

def inhand(inhand_obj:item):
  return holds_rh(char, inhand_obj) or holds_lh(char, inhand_obj)

def standing(char: character):
  return not sitting(char) and not lying(char)

def has_a_free_hand():
  symbol l=exists item1: item : holds_lh(char, item1)
  symbol r=exists item2: item : holds_rh(char, item2)
  return not l or not r



behavior put(inhand_obj: item, obj: item):
  body:
    assert surfaces(obj) or is_room(obj) or recipient(obj) or containers(obj) or can_open(obj) or eatable(obj)
    achieve inhand(inhand_obj)
    if can_open(obj) and closed(obj):
      achieve open(obj)
    achieve close_char(char, obj)
    put_executor(inhand_obj, obj)

  eff:
    holds_rh[char, inhand_obj] = False
    holds_lh[char, inhand_obj] = False
    if surfaces(obj):
      on[inhand_obj, obj] = True
    if is_room(obj) or recipient(obj) or containers(obj) or can_open(obj):
      inside[inhand_obj, obj] = True
    close[inhand_obj, obj] = True
    close[obj, inhand_obj] = True
    foreach inter in (findall x: item: close(x, obj)):
      close[inter, inhand_obj] = True
      close[inhand_obj, inter] = True

behavior empty_a_hand():
  goal: has_a_free_hand()
  body:
    assert not has_a_free_hand()
    bind surf:item where:
      surfaces(surf)
    bind give_up_obj:item where:
      inhand(give_up_obj)
    put(give_up_obj, surf)

behavior stand():
  goal: standing(char)
  body:
    assert sitting(char) or lying(char)
    standup_executor(char)
  eff:
    sitting[char] = False
    lying[char] = False

behavior sit():
  goal: sitting(char)
  body:
    assert not sitting(char)
    bind seat:item where:
      sittable(seat)
    achieve close_char(char, seat)
    sit_executor(seat)
  eff:
    sitting[char] = True
    on_char[char, seat] = True
    lying[char] = False

behavior lie():
  goal: lying(char)
  body:
    assert not lying(char)
    bind bed:item where:
      lieable(bed)
    achieve close_char(char, bed)
    lie_executor(bed)
  eff:
    lying[char] = True
    sitting[char] = False
    on_char[char, bed] = True

def obj_inside_or_on(obj1: item, obj2: item):
  return inside(obj1, obj2) or on(obj2, obj1)

behavior walk(obj: item):
  goal: close_char(char, obj)
  body:
    achieve standing(char)
    walk_executor(obj)
    let inhand_objects=findall o: item where: inhand(o)

  eff:
    # foreach icf:item:
    #   inside_char[char,icf]= False
    #   close_char[char, icf]= False
    #   facing_char[char, icf]= False
    #   foreach o in inhand_objects:
    #     inside[o, icf] = False
    #     close[o, icf] = False
    #     close[icf, o] = False
    #     facing[o, icf] = False
    #     facing[icf, o] = False

    #   if obj_inside_or_on(obj, icf):
    #     close_char[char, icf] = True
    #     foreach o in inhand_objects:
    #       close[o, icf] = True
    #       close[icf, o] = True

    inside_char[char, :] = False
    close_char[char, :] = False
    facing_char[char, :] = False
    foreach o in inhand_objects:
      inside[o, :]= False
      close[o, :] = False
      close[:, o] = False

    foreach icf in (findall t:item: obj_inside_or_on(obj, t)):
      close_char[char, icf] = True
      foreach o in inhand_objects:
        close[o, icf] = True
        close[icf, o] = True

    close_char[char,obj] = True
    foreach o in inhand_objects:
      close[o, obj] = True
      close[obj, o] = True

behavior find(obj:item):
  goal: facing_char(char, obj) and close_char(char, obj)
  body:
    if on_body(obj, char):
      find_executor(obj)
    else:
      achieve close_char(char, obj)
      find_executor(obj)
  eff:
    foreach o in (findall t:item: facing_char(char, t)):
      facing_char[char, o] = False
    facing_char[char, obj] = True

behavior turnto(obj:item):
  goal: facing_char(char, obj)
  body:
    turnto_executor(obj)
  eff:
    foreach o in (findall t:item: facing_char(char, t)):
      facing_char[char, o] = False
    facing_char[char, obj] = True

behavior switch_off(obj: item):
  goal: is_off(obj)
  body:
    assert has_switch(obj)
    assert is_on(obj)
    achieve has_a_free_hand()
    achieve close_char(char, obj)
    switchoff_executor(obj)
  eff:
    is_off[obj] = True
    is_on[obj] = False

behavior switch_on(obj: item):
  goal: is_on(obj)
  body:
    assert has_switch(obj)
    achieve has_a_free_hand()
    if has_plug(obj):
      achieve plugged(obj)
    if can_open(obj):
      achieve closed(obj)
    achieve close_char(char, obj)
    switchon_executor(obj)
  eff:
    is_off[obj] = False
    is_on[obj] = True

behavior put_close(inhand_obj: item, obj: item):
  goal: close(inhand_obj, obj)
  body:
    put(inhand_obj, obj)

behavior put_on(inhand_obj: item, obj: item):
  goal: on(inhand_obj, obj)
  body:
    put(inhand_obj, obj)


behavior put_inside(inhand_obj: item, obj: item):
  goal: inside(inhand_obj, obj)
  body:
    put(inhand_obj, obj)

behavior grab(obj: item):
  goal: inhand(obj)
  body:
    assert grabbable(obj) or is_water(obj)
    achieve has_a_free_hand()
    foreach obj2:item:
      if inside(obj,obj2):
        if not is_room(obj2):
          assert can_open(obj2) or recipient(obj2) or eatable(obj2)
          if can_open(obj2):
            achieve open(obj2)
    achieve close_char(char, obj)
    grab_executor(obj)
  eff:
    on[obj, :] = False
    on[:, obj] = False
    inside[obj, :] = False
    inside[:, obj] = False
    close[obj, :] = False
    close[:, obj] = False
    if exists item1: item : holds_lh(char, item1):
      holds_rh[char, obj] = True
    else:
      holds_lh[char, obj] = True
    close_char[char,obj]=True

behavior wash(obj: item):
  goal: clean(obj)
  body:
    achieve has_a_free_hand()
    achieve close_char(char, obj)
    wash_executor(obj)
  eff:
    dirty[obj] = False
    clean[obj] = True

behavior open(obj: item):
  goal: open(obj)
  body:
    assert can_open(obj)
    assert closed(obj)
    achieve has_a_free_hand()
    if has_switch(obj):
      achieve is_off(obj)
    achieve close_char(char, obj)
    open_executor(obj)
  eff:
    open[obj] = True
    closed[obj] = False

behavior closes(obj: item):
  goal: closed(obj)
  body:
    assert can_open(obj)
    assert open(obj)
    achieve has_a_free_hand()
    achieve close_char(char, obj)
    close_executor(obj)
  eff:
    open[obj] = False
    closed[obj] = True

def pour_target(obj: item):
  return is_hands_both(obj) or is_sponge(obj) or is_face(obj)

behavior pour(obj: item, target: item):
  goal: inside(obj, target)
  body:

    assert pourable(obj) or drinkable(obj)
    assert recipient(target) or pour_target(obj)
    achieve inhand(obj)
    achieve close_char(char, target)
    pour_executor(obj, target)
  eff:
    inside[obj, target] = True
    if is_water(obj):
      holds_lh[char, obj] = False
      holds_rh[char, obj] = False

behavior plugin(object:item):
  goal: plugged(object)
  body:
    assert has_plug(object)
    achieve has_a_free_hand()
    achieve close_char(char, object)
    plugin_executor(object)
  eff:
    plugged[object] = True
    unplugged[object] = False

behavior plugout(object:item):
  goal: unplugged(object)
  body:
    assert has_plug(object)
    achieve has_a_free_hand()
    if has_switch(object):
      achieve is_off(object)
    achieve close_char(char, object)
    plugout_executor(object)
  eff:
    plugged[object] = False
    unplugged[object] = True

behavior cut(object:item):
  goal: cut(object)
  body:
    assert cuttable(object) or eatable(object)
    achieve has_a_free_hand()
    symbol has_knife=exists knife:item: is_knife(knife) and inhand(knife)
    if not has_knife:
      bind new_knife:item where:
        is_knife(new_knife)
      achieve inhand(new_knife)
    achieve close_char(char, object)
    cut_executor(object)
  eff:
    cut[object] = True

behavior eat(object:item):
  body:
    assert eatable(object)
    eat_executor(object)


behavior sleep():
  goal: sleeping(char)
  body:
    symbol has_lieable_place=exists item1:item: lieable(item1)
    symbol has_sittable_place=exists item2:item: sittable(item2)
    assert has_lieable_place or has_sittable_place
    if has_lieable_place:
      lie()
    else:
      sit()
  eff:
    sleeping[char] = True

behavior wake_up():
  goal: not sleeping(char)
  body:
    assert sleeping(char)
    stand()
  eff:
    sleeping[char] = False

behavior wipe(obj:item):
  goal: clean(obj)
  body:
    symbol has_cleaning_solution=exists item1:item: is_towel(item1) or is_rag(item1) or is_sponge(item1) or is_paper_towel(item1) or is_cloth_napkin(item1) or is_duster(item1) or is_cleaning_solution(item1)
    if not has_cleaning_solution:
      bind cleaning_tool:item where:
        is_towel(cleaning_tool) or is_rag(cleaning_tool) or is_sponge(cleaning_tool) or is_paper_towel(cleaning_tool) or is_cloth_napkin(cleaning_tool) or is_duster(cleaning_tool) or is_cleaning_solution(cleaning_tool)
      achieve inhand(cleaning_tool)
    achieve close_char(char, obj)
    wipe_executor(obj)
  eff:
    dirty[obj] = False
    clean[obj] = True

behavior put_on_body(inhand_obj: item):
  goal: on_body(inhand_obj, char)
  body:
    assert clothes(inhand_obj)
    achieve inhand(inhand_obj)
    puton_executor(inhand_obj)
  eff:
    on_body[inhand_obj, char] = True

behavior put_off_body(clo: item):
  goal: not on_body(clo, char)
  body:
    assert clothes(clo)
    putoff_executor(clo)
  eff:
    on_body[clo, char] = False

behavior read(material:item):
  body:
    assert readable(material)
    achieve inhand(material)
    read_executor(material)

behavior touch(obj:item):
  body:
    foreach obj2:item:
      if inside(obj,obj2):
        if not is_room(obj2):
          assert can_open(obj2) or recipient(obj2) or eatable(obj2)
          if can_open(obj2):
            achieve open(obj2)
    achieve close_char(char, obj)
    touch_executor(obj)

behavior type(obj:item):
  body:
    assert is_keyboard(obj) or has_switch(obj)
    achieve close_char(char, obj)
    type_executor(obj)

behavior watch(obj:item):
  body:
    assert lookable(obj)
    achieve facing_char(char, obj)

behavior drink(obj: item):
  body:
    assert drinkable(obj) or recipient(obj)
    achieve inhand(obj)
    drink_executor(obj)

behavior look_at(obj:item):
  body:
    achieve facing_char(char, obj)
    lookat_executor(obj)

behavior greet(person:item):
  body:
    assert person(person)
    greet_executor(person)

behavior move(obj:item):
  body:
    assert movable(obj) or is_button(obj) or is_chair(obj) or is_curtain(obj)
    achieve has_a_free_hand()
    achieve close_char(char, obj)
    move_executor(obj)

behavior squeeze(obj:item):
  body:
    assert is_cleaning_solution(obj) or is_tooth_paste(obj) or is_shampoo(obj) or is_sponge(obj) or clothes(obj)
    achieve has_a_free_hand()
    achieve close_char(char, obj)
