problem "agent-problem"
domain "virtualhome_partial.cdl"

#!pragma planner_is_goal_serializable=False
#!pragma planner_is_goal_ordered=True
#!pragma planner_always_commit_skeleton=True

objects:
#objects
  clothes_pants_2157:item
  clothes_shirt_2158:item
  clothes_socks_2159:item
  clothes_skirt_2160:item
  iron_2161:item
  basket_for_clothes_2078:item
  washing_machine_2079:item
  food_steak_2080:item
  food_apple_2081:item
  food_bacon_2082:item
  food_banana_2083:item
  food_bread_2084:item
  food_cake_2085:item
  food_carrot_2086:item
  food_cereal_2087:item
  food_cheese_2088:item
  food_chicken_2089:item
  food_dessert_2090:item
  food_donut_2091:item
  food_egg_2092:item
  food_fish_2093:item
  food_food_2094:item
  food_fruit_2095:item
  food_hamburger_2096:item
  food_ice_cream_2097:item
  food_jam_2098:item
  food_kiwi_2099:item
  food_lemon_2100:item
  food_noodles_2101:item
  food_oatmeal_2102:item
  food_orange_2103:item
  food_onion_2104:item
  food_peanut_butter_2105:item
  food_pizza_2106:item
  food_potato_2107:item
  food_rice_2108:item
  food_salt_2109:item
  food_snack_2110:item
  food_sugar_2111:item
  food_turkey_2112:item
  food_vegetable_2113:item
  dry_pasta_2114:item
  milk_2115:item
  clothes_dress_2116:item
  clothes_hat_2117:item
  clothes_gloves_2118:item
  clothes_jacket_2119:item
  clothes_scarf_2120:item
  clothes_underwear_2121:item
  knife_2122:item
  cutting_board_2123:item
  remote_control_2124:item
  soap_2125:item
  soap_2126:item
  towel_2128:item
  cd_player_2129:item
  dvd_player_2130:item
  headset_2131:item
  cup_2132:item
  cup_2133:item
  cup_2134:item
  stove_2135:item
  book_2136:item
  book_2137:item
  pot_2138:item
  vacuum_cleaner_2139:item
  bowl_2140:item
  bowl_2141:item
  bowl_2142:item
  cleaning_solution_2143:item
  ironing_board_2144:item
  cd_2145:item
  headset_2146:item
  phone_2147:item
  sauce_2148:item
  oil_2149:item
  fork_2150:item
  fork_2151:item
  plate_2152:item
  spectacles_2153:item
  fryingpan_2154:item
  detergent_2155:item
  window_2156:item
  bathroom_1:item
  wall_2:item
  wall_3:item
  wall_4:item
  wall_5:item
  ceiling_6:item
  ceiling_7:item
  ceiling_8:item
  ceiling_9:item
  floor_10:item
  floor_11:item
  floor_12:item
  floor_13:item
  floor_14:item
  toilet_15:item
  shower_16:item
  bathroom_cabinet_17:item
  bathroom_counter_18:item
  sink_19:item
  faucet_20:item
  shower_21:item
  curtain_22:item
  mat_32:item
  drawing_33:item
  walllamp_34:item
  ceilinglamp_35:item
  walllamp_36:item
  doorjamb_37:item
  door_38:item
  light_39:item
  dining_room_41:item
  floor_42:item
  floor_43:item
  floor_44:item
  floor_45:item
  floor_46:item
  floor_47:item
  floor_48:item
  floor_49:item
  floor_50:item
  floor_51:item
  ceiling_52:item
  ceiling_53:item
  ceiling_54:item
  ceiling_55:item
  ceiling_56:item
  ceiling_57:item
  ceiling_58:item
  ceiling_59:item
  ceiling_60:item
  door_61:item
  door_62:item
  wall_63:item
  wall_64:item
  wall_65:item
  wall_66:item
  wall_67:item
  wall_68:item
  wall_69:item
  wall_70:item
  phone_71:item
  powersocket_72:item
  light_73:item
  knifeblock_76:item
  pot_78:item
  trashcan_99:item
  mat_102:item
  pillow_103:item
  pillow_104:item
  pillow_105:item
  pillow_106:item
  pillow_107:item
  pillow_108:item
  drawing_110:item
  drawing_111:item
  bench_113:item
  table_114:item
  bench_115:item
  tvstand_116:item
  cupboard_117:item
  cupboard_118:item
  kitchen_counter_119:item
  sink_120:item
  faucet_121:item
  kitchen_counter_122:item
  kitchen_counter_123:item
  bookshelf_124:item
  stovefan_125:item
  fridge_126:item
  oven_127:item
  tray_128:item
  dishwasher_129:item
  coffe_maker_130:item
  toaster_132:item
  microwave_135:item
  ceilinglamp_137:item
  ceilinglamp_138:item
  walllamp_139:item
  walllamp_140:item
  walllamp_141:item
  bedroom_162:item
  floor_163:item
  floor_164:item
  floor_165:item
  floor_166:item
  floor_167:item
  floor_168:item
  floor_169:item
  floor_170:item
  floor_171:item
  floor_172:item
  wall_173:item
  wall_174:item
  wall_175:item
  wall_176:item
  wall_177:item
  wall_178:item
  wall_179:item
  wall_180:item
  ceiling_181:item
  ceiling_182:item
  ceiling_183:item
  ceiling_184:item
  ceiling_185:item
  ceiling_186:item
  ceiling_187:item
  ceiling_188:item
  ceiling_189:item
  doorjamb_190:item
  window_191:item
  nightstand_192:item
  desk_193:item
  chair_194:item
  nightstand_195:item
  bookshelf_196:item
  bed_197:item
  couch_198:item
  table_199:item
  filing_cabinet_200:item
  drawing_201:item
  drawing_202:item
  mat_203:item
  curtain_204:item
  curtain_205:item
  curtain_206:item
  pillow_207:item
  pillow_208:item
  computer_209:item
  cpuscreen_210:item
  keyboard_211:item
  light_212:item
  mouse_213:item
  mousepad_214:item
  photoframe_219:item
  ceilinglamp_237:item
  tablelamp_238:item
  tablelamp_239:item
  home_office_241:item
  wall_242:item
  wall_243:item
  wall_244:item
  wall_245:item
  wall_246:item
  wall_247:item
  wall_248:item
  wall_249:item
  ceiling_250:item
  ceiling_251:item
  ceiling_252:item
  ceiling_253:item
  ceiling_254:item
  ceiling_255:item
  ceiling_256:item
  ceiling_257:item
  ceiling_258:item
  floor_259:item
  floor_260:item
  floor_261:item
  floor_262:item
  floor_263:item
  floor_264:item
  floor_265:item
  floor_266:item
  floor_267:item
  floor_268:item
  couch_269:item
  table_270:item
  chair_271:item
  desk_272:item
  tvstand_273:item
  dresser_274:item
  bookshelf_275:item
  computer_276:item
  cpuscreen_277:item
  keyboard_278:item
  mousepad_279:item
  mouse_280:item
  television_281:item
  powersocket_282:item
  light_283:item
  mat_284:item
  orchid_285:item
  pillow_286:item
  pillow_287:item
  drawing_288:item
  curtain_289:item
  curtain_290:item
  curtain_291:item
  hanger_292:item
  hanger_293:item
  hanger_294:item
  ceilinglamp_303:item
  walllamp_304:item
  walllamp_305:item
  walllamp_306:item
  walllamp_307:item
  doorjamb_308:item
  doorjamb_309:item
  window_310:item
  food_food_1000:item
  wooden_spoon_2000:item
  food_food_2001:item
  brush_2002:item
  chair_2003:item
  lighter_2004:item
  table_cloth_2005:item
  piano_bench_2006:item
  food_butter_2007:item
  diary_2008:item
  food_onion_2009:item
  soap_2010:item
  detergent_2011:item
  measuring_cup_2012:item
  oil_2013:item
  pencil_2014:item
  food_carrot_2015:item
  phone_2016:item
  phone_2017:item
  envelope_2018:item
  shampoo_2019:item
  pencil_2020:item
  food_food_2021:item
  stamp_2022:item
  tea_bag_2023:item
  ice_2024:item
  rag_2025:item
  check_2026:item
  food_orange_2027:item
  instrument_guitar_2028:item
  phone_2029:item
  cd_2030:item
  scrabble_2031:item
  shoes_2033:item
  laser_pointer_2034:item
  knife_2035:item
  clothes_pants_2036:item
  knife_2037:item
  box_2038:item
  lighter_2039:item
  pot_2040:item
  food_salt_2041:item
  after_shave_2042:item
  stamp_2043:item
  shoe_rack_2044:item
  glue_2045:item
  food_food_2046:item
  homework_2047:item
  food_onion_2048:item
  cup_2049:item
  stereo_2050:item
  after_shave_2051:item
  rag_2052:item
  coffee_filter_2053:item
  food_kiwi_2054:item
  envelope_2055:item
  toy_2056:item
  blow_dryer_2057:item
  check_2058:item
  tooth_paste_2059:item
  novel_2060:item
  food_orange_2061:item
  piano_bench_2062:item
  after_shave_2063:item
  food_food_2064:item
  coffee_filter_2065:item
  tea_2066:item
  piano_bench_2067:item
  tray_2068:item
  cat_2069:item
  chessboard_2070:item
  check_2071:item
  food_cheese_2072:item
  food_food_2073:item
  food_food_2074:item
  check_2075:item
  toilet_paper_2076:item
  food_peanut_butter_2077:item
#object_end

init:
    #categories
    is_pants[clothes_pants_2157]=True
    is_clothes_pants[clothes_pants_2157]=True
    is_clothes_shirt[clothes_shirt_2158]=True
    is_shirt[clothes_shirt_2158]=True
    is_clothes_socks[clothes_socks_2159]=True
    is_clothes_skirt[clothes_skirt_2160]=True
    is_iron[iron_2161]=True
    is_clothes_pile[basket_for_clothes_2078]=True
    is_basket_for_clothes[basket_for_clothes_2078]=True
    is_washing_machine[washing_machine_2079]=True
    is_food_steak[food_steak_2080]=True
    is_food_apple[food_apple_2081]=True
    is_apple[food_apple_2081]=True
    is_food_bacon[food_bacon_2082]=True
    is_food_banana[food_banana_2083]=True
    is_banana[food_banana_2083]=True
    is_bread_slice[food_bread_2084]=True
    is_bread[food_bread_2084]=True
    is_food_bread[food_bread_2084]=True
    is_food_cake[food_cake_2085]=True
    is_food_carrot[food_carrot_2086]=True
    is_carrot[food_carrot_2086]=True
    is_cereal[food_cereal_2087]=True
    is_food_cereal[food_cereal_2087]=True
    is_food_cheese[food_cheese_2088]=True
    is_food_chicken[food_chicken_2089]=True
    is_chicken[food_chicken_2089]=True
    is_pie[food_dessert_2090]=True
    is_creamybuns[food_dessert_2090]=True
    is_pancake[food_dessert_2090]=True
    is_cupcake[food_dessert_2090]=True
    is_watermelon[food_dessert_2090]=True
    is_milkshake[food_dessert_2090]=True
    is_poundcake[food_dessert_2090]=True
    is_sundae[food_dessert_2090]=True
    is_pudding[food_dessert_2090]=True
    is_food_dessert[food_dessert_2090]=True
    is_food_donut[food_donut_2091]=True
    is_food_egg[food_egg_2092]=True
    is_food_fish[food_fish_2093]=True
    is_salmon[food_fish_2093]=True
    is_creamybuns[food_food_2094]=True
    is_cutlets[food_food_2094]=True
    is_salmon[food_food_2094]=True
    is_pear[food_food_2094]=True
    is_chicken[food_food_2094]=True
    is_plum[food_food_2094]=True
    is_orange[food_food_2094]=True
    is_cereal[food_food_2094]=True
    is_banana[food_food_2094]=True
    is_bell_pepper[food_food_2094]=True
    is_apple[food_food_2094]=True
    is_whippedcream[food_food_2094]=True
    is_chinesefood[food_food_2094]=True
    is_food_food[food_food_2094]=True
    is_tomato[food_food_2094]=True
    is_bananas[food_food_2094]=True
    is_chocolatesyrup[food_food_2094]=True
    is_potato[food_food_2094]=True
    is_bellpepper[food_food_2094]=True
    is_crackers[food_food_2094]=True
    is_cucumber[food_food_2094]=True
    is_plum[food_fruit_2095]=True
    is_food_fruit[food_fruit_2095]=True
    is_orange[food_fruit_2095]=True
    is_banana[food_fruit_2095]=True
    is_watermelon[food_fruit_2095]=True
    is_apple[food_fruit_2095]=True
    is_pear[food_fruit_2095]=True
    is_mincedmeat[food_hamburger_2096]=True
    is_food_hamburger[food_hamburger_2096]=True
    is_food_ice_cream[food_ice_cream_2097]=True
    is_food_jam[food_jam_2098]=True
    is_food_kiwi[food_kiwi_2099]=True
    is_food_lemon[food_lemon_2100]=True
    is_lemon[food_lemon_2100]=True
    is_food_noodles[food_noodles_2101]=True
    is_food_oatmeal[food_oatmeal_2102]=True
    is_cereal[food_oatmeal_2102]=True
    is_food_orange[food_orange_2103]=True
    is_food_onion[food_onion_2104]=True
    is_food_peanut_butter[food_peanut_butter_2105]=True
    is_food_pizza[food_pizza_2106]=True
    is_potato[food_potato_2107]=True
    is_food_potato[food_potato_2107]=True
    is_food_rice[food_rice_2108]=True
    is_condiment_shaker[food_salt_2109]=True
    is_food_salt[food_salt_2109]=True
    is_salt_crackers[food_snack_2110]=True
    is_chips[food_snack_2110]=True
    is_cupcake[food_snack_2110]=True
    is_candybar[food_snack_2110]=True
    is_banana[food_snack_2110]=True
    is_crackers[food_snack_2110]=True
    is_food_snack[food_snack_2110]=True
    is_poundcake[food_snack_2110]=True
    is_apple[food_snack_2110]=True
    is_condiment_shaker[food_sugar_2111]=True
    is_food_sugar[food_sugar_2111]=True
    is_food_turkey[food_turkey_2112]=True
    is_chicken[food_turkey_2112]=True
    is_food_vegetable[food_vegetable_2113]=True
    is_salad[food_vegetable_2113]=True
    is_potato[food_vegetable_2113]=True
    is_carrot[food_vegetable_2113]=True
    is_tomato[food_vegetable_2113]=True
    is_cucumber[food_vegetable_2113]=True
    is_dry_pasta[dry_pasta_2114]=True
    is_milk[milk_2115]=True
    is_clothes_dress[clothes_dress_2116]=True
    is_clothes_hat[clothes_hat_2117]=True
    is_clothes_gloves[clothes_gloves_2118]=True
    is_clothes_jacket[clothes_jacket_2119]=True
    is_clothes_scarf[clothes_scarf_2120]=True
    is_clothes_underwear[clothes_underwear_2121]=True
    is_chefknife[knife_2122]=True
    is_cutlery_knife[knife_2122]=True
    is_knife[knife_2122]=True
    is_cutting_board[cutting_board_2123]=True
    is_remote_control[remote_control_2124]=True
    is_controller[remote_control_2124]=True
    is_soap[soap_2125]=True
    is_barsoap[soap_2125]=True
    is_soap[soap_2126]=True
    is_barsoap[soap_2126]=True
    is_towel[towel_2128]=True
    is_radio[cd_player_2129]=True
    is_cd_player[cd_player_2129]=True
    is_dvd_player[dvd_player_2130]=True
    is_headset[headset_2131]=True
    is_wineglass[cup_2132]=True
    is_cup[cup_2132]=True
    is_waterglass[cup_2132]=True
    is_mug[cup_2132]=True
    is_wineglass[cup_2133]=True
    is_cup[cup_2133]=True
    is_waterglass[cup_2133]=True
    is_mug[cup_2133]=True
    is_wineglass[cup_2134]=True
    is_cup[cup_2134]=True
    is_waterglass[cup_2134]=True
    is_mug[cup_2134]=True
    is_oven[stove_2135]=True
    is_stove[stove_2135]=True
    is_book[book_2136]=True
    is_textbook[book_2136]=True
    is_novel[book_2136]=True
    is_book[book_2137]=True
    is_textbook[book_2137]=True
    is_novel[book_2137]=True
    is_pot[pot_2138]=True
    is_vacuum_cleaner[vacuum_cleaner_2139]=True
    is_bowl[bowl_2140]=True
    is_dish_bowl[bowl_2140]=True
    is_bowl[bowl_2141]=True
    is_dish_bowl[bowl_2141]=True
    is_bowl[bowl_2142]=True
    is_dish_bowl[bowl_2142]=True
    is_cleaning_solution[cleaning_solution_2143]=True
    is_dishwashingliquid[cleaning_solution_2143]=True
    is_ironing_board[ironing_board_2144]=True
    is_cd[cd_2145]=True
    is_headset[headset_2146]=True
    is_wall_phone[phone_2147]=True
    is_phone[phone_2147]=True
    is_cellphone[phone_2147]=True
    is_sauce[sauce_2148]=True
    is_condiment_bottle[sauce_2148]=True
    is_oil[oil_2149]=True
    is_condiment_bottle[oil_2149]=True
    is_fork[fork_2150]=True
    is_cutlery_fork[fork_2150]=True
    is_fork[fork_2151]=True
    is_cutlery_fork[fork_2151]=True
    is_plate[plate_2152]=True
    is_glasses[spectacles_2153]=True
    is_spectacles[spectacles_2153]=True
    is_fryingpan[fryingpan_2154]=True
    is_dishwashingliquid[detergent_2155]=True
    is_detergent[detergent_2155]=True
    is_window[window_2156]=True
    is_bathroom[bathroom_1]=True
    is_wall[wall_2]=True
    is_wall[wall_3]=True
    is_wall[wall_4]=True
    is_wall[wall_5]=True
    is_ceiling[ceiling_6]=True
    is_ceiling[ceiling_7]=True
    is_ceiling[ceiling_8]=True
    is_ceiling[ceiling_9]=True
    is_floor[floor_10]=True
    is_floor[floor_11]=True
    is_floor[floor_12]=True
    is_floor[floor_13]=True
    is_floor[floor_14]=True
    is_toilet[toilet_15]=True
    is_stall[shower_16]=True
    is_shower[shower_16]=True
    is_bathroom_cabinet[bathroom_cabinet_17]=True
    is_bathroom_counter[bathroom_counter_18]=True
    is_sink[sink_19]=True
    is_faucet[faucet_20]=True
    is_stall[shower_21]=True
    is_shower[shower_21]=True
    is_curtains[curtain_22]=True
    is_curtain[curtain_22]=True
    is_rug[mat_32]=True
    is_mat[mat_32]=True
    is_drawing[drawing_33]=True
    is_wallpictureframe[drawing_33]=True
    is_walllamp[walllamp_34]=True
    is_ceilinglamp[ceilinglamp_35]=True
    is_walllamp[walllamp_36]=True
    is_doorjamb[doorjamb_37]=True
    is_door[door_38]=True
    is_light_switch[light_39]=True
    is_lightswitch[light_39]=True
    is_light[light_39]=True
    is_kitchen[dining_room_41]=True
    is_dining_room[dining_room_41]=True
    is_floor[floor_42]=True
    is_floor[floor_43]=True
    is_floor[floor_44]=True
    is_floor[floor_45]=True
    is_floor[floor_46]=True
    is_floor[floor_47]=True
    is_floor[floor_48]=True
    is_floor[floor_49]=True
    is_floor[floor_50]=True
    is_floor[floor_51]=True
    is_ceiling[ceiling_52]=True
    is_ceiling[ceiling_53]=True
    is_ceiling[ceiling_54]=True
    is_ceiling[ceiling_55]=True
    is_ceiling[ceiling_56]=True
    is_ceiling[ceiling_57]=True
    is_ceiling[ceiling_58]=True
    is_ceiling[ceiling_59]=True
    is_ceiling[ceiling_60]=True
    is_door[door_61]=True
    is_door[door_62]=True
    is_wall[wall_63]=True
    is_wall[wall_64]=True
    is_wall[wall_65]=True
    is_wall[wall_66]=True
    is_wall[wall_67]=True
    is_wall[wall_68]=True
    is_wall[wall_69]=True
    is_wall[wall_70]=True
    is_wall_phone[phone_71]=True
    is_phone[phone_71]=True
    is_cellphone[phone_71]=True
    is_powersocket[powersocket_72]=True
    is_light_switch[light_73]=True
    is_lightswitch[light_73]=True
    is_light[light_73]=True
    is_knifeblock[knifeblock_76]=True
    is_pot[pot_78]=True
    is_trashcan[trashcan_99]=True
    is_garbage_can[trashcan_99]=True
    is_rug[mat_102]=True
    is_mat[mat_102]=True
    is_pillow[pillow_103]=True
    is_pillow[pillow_104]=True
    is_pillow[pillow_105]=True
    is_pillow[pillow_106]=True
    is_pillow[pillow_107]=True
    is_pillow[pillow_108]=True
    is_drawing[drawing_110]=True
    is_wallpictureframe[drawing_110]=True
    is_drawing[drawing_111]=True
    is_wallpictureframe[drawing_111]=True
    is_bench[bench_113]=True
    is_coffee_table[table_114]=True
    is_diningtable[table_114]=True
    is_table[table_114]=True
    is_kitchen_table[table_114]=True
    is_bench[bench_115]=True
    is_tvstand[tvstand_116]=True
    is_cupboard[cupboard_117]=True
    is_kitchen_cabinets[cupboard_117]=True
    is_cupboard[cupboard_118]=True
    is_kitchen_cabinets[cupboard_118]=True
    is_kitchen_counter[kitchen_counter_119]=True
    is_sink[sink_120]=True
    is_faucet[faucet_121]=True
    is_kitchen_counter[kitchen_counter_122]=True
    is_kitchen_counter[kitchen_counter_123]=True
    is_bookshelf[bookshelf_124]=True
    is_stovefan[stovefan_125]=True
    is_freezer[fridge_126]=True
    is_fridge[fridge_126]=True
    is_oven[oven_127]=True
    is_stove[oven_127]=True
    is_oventray[tray_128]=True
    is_tray[tray_128]=True
    is_dishwasher[dishwasher_129]=True
    is_coffe_maker[coffe_maker_130]=True
    is_coffeemaker[coffe_maker_130]=True
    is_toaster[toaster_132]=True
    is_microwave[microwave_135]=True
    is_ceilinglamp[ceilinglamp_137]=True
    is_ceilinglamp[ceilinglamp_138]=True
    is_walllamp[walllamp_139]=True
    is_walllamp[walllamp_140]=True
    is_walllamp[walllamp_141]=True
    is_bedroom[bedroom_162]=True
    is_floor[floor_163]=True
    is_floor[floor_164]=True
    is_floor[floor_165]=True
    is_floor[floor_166]=True
    is_floor[floor_167]=True
    is_floor[floor_168]=True
    is_floor[floor_169]=True
    is_floor[floor_170]=True
    is_floor[floor_171]=True
    is_floor[floor_172]=True
    is_wall[wall_173]=True
    is_wall[wall_174]=True
    is_wall[wall_175]=True
    is_wall[wall_176]=True
    is_wall[wall_177]=True
    is_wall[wall_178]=True
    is_wall[wall_179]=True
    is_wall[wall_180]=True
    is_ceiling[ceiling_181]=True
    is_ceiling[ceiling_182]=True
    is_ceiling[ceiling_183]=True
    is_ceiling[ceiling_184]=True
    is_ceiling[ceiling_185]=True
    is_ceiling[ceiling_186]=True
    is_ceiling[ceiling_187]=True
    is_ceiling[ceiling_188]=True
    is_ceiling[ceiling_189]=True
    is_doorjamb[doorjamb_190]=True
    is_window[window_191]=True
    is_nightstand[nightstand_192]=True
    is_cpu_table[desk_193]=True
    is_desk[desk_193]=True
    is_chair[chair_194]=True
    is_nightstand[nightstand_195]=True
    is_bookshelf[bookshelf_196]=True
    is_bed[bed_197]=True
    is_couch[couch_198]=True
    is_sofa[couch_198]=True
    is_coffee_table[table_199]=True
    is_diningtable[table_199]=True
    is_table[table_199]=True
    is_kitchen_table[table_199]=True
    is_filing_cabinet[filing_cabinet_200]=True
    is_cabinet[filing_cabinet_200]=True
    is_drawing[drawing_201]=True
    is_wallpictureframe[drawing_201]=True
    is_drawing[drawing_202]=True
    is_wallpictureframe[drawing_202]=True
    is_rug[mat_203]=True
    is_mat[mat_203]=True
    is_curtains[curtain_204]=True
    is_curtain[curtain_204]=True
    is_curtains[curtain_205]=True
    is_curtain[curtain_205]=True
    is_curtains[curtain_206]=True
    is_curtain[curtain_206]=True
    is_pillow[pillow_207]=True
    is_pillow[pillow_208]=True
    is_cpu_case[computer_209]=True
    is_computer[computer_209]=True
    is_pc[computer_209]=True
    is_cpuscreen[cpuscreen_210]=True
    is_keyboard[keyboard_211]=True
    is_light_switch[light_212]=True
    is_lightswitch[light_212]=True
    is_light[light_212]=True
    is_mouse[mouse_213]=True
    is_mouse_mat[mousepad_214]=True
    is_mousemat[mousepad_214]=True
    is_mousepad[mousepad_214]=True
    is_photoframe[photoframe_219]=True
    is_ceilinglamp[ceilinglamp_237]=True
    is_tablelamp[tablelamp_238]=True
    is_tablelamp[tablelamp_239]=True
    is_livingroom[home_office_241]=True
    is_home_office[home_office_241]=True
    is_wall[wall_242]=True
    is_wall[wall_243]=True
    is_wall[wall_244]=True
    is_wall[wall_245]=True
    is_wall[wall_246]=True
    is_wall[wall_247]=True
    is_wall[wall_248]=True
    is_wall[wall_249]=True
    is_ceiling[ceiling_250]=True
    is_ceiling[ceiling_251]=True
    is_ceiling[ceiling_252]=True
    is_ceiling[ceiling_253]=True
    is_ceiling[ceiling_254]=True
    is_ceiling[ceiling_255]=True
    is_ceiling[ceiling_256]=True
    is_ceiling[ceiling_257]=True
    is_ceiling[ceiling_258]=True
    is_floor[floor_259]=True
    is_floor[floor_260]=True
    is_floor[floor_261]=True
    is_floor[floor_262]=True
    is_floor[floor_263]=True
    is_floor[floor_264]=True
    is_floor[floor_265]=True
    is_floor[floor_266]=True
    is_floor[floor_267]=True
    is_floor[floor_268]=True
    is_couch[couch_269]=True
    is_sofa[couch_269]=True
    is_coffee_table[table_270]=True
    is_diningtable[table_270]=True
    is_table[table_270]=True
    is_kitchen_table[table_270]=True
    is_chair[chair_271]=True
    is_cpu_table[desk_272]=True
    is_desk[desk_272]=True
    is_tvstand[tvstand_273]=True
    is_closet[dresser_274]=True
    is_dresser[dresser_274]=True
    is_bookshelf[bookshelf_275]=True
    is_cpu_case[computer_276]=True
    is_computer[computer_276]=True
    is_pc[computer_276]=True
    is_cpuscreen[cpuscreen_277]=True
    is_keyboard[keyboard_278]=True
    is_mouse_mat[mousepad_279]=True
    is_mousemat[mousepad_279]=True
    is_mousepad[mousepad_279]=True
    is_mouse[mouse_280]=True
    is_walltv[television_281]=True
    is_television[television_281]=True
    is_tv[television_281]=True
    is_powersocket[powersocket_282]=True
    is_light_switch[light_283]=True
    is_lightswitch[light_283]=True
    is_light[light_283]=True
    is_rug[mat_284]=True
    is_mat[mat_284]=True
    is_orchid[orchid_285]=True
    is_pillow[pillow_286]=True
    is_pillow[pillow_287]=True
    is_drawing[drawing_288]=True
    is_wallpictureframe[drawing_288]=True
    is_curtains[curtain_289]=True
    is_curtain[curtain_289]=True
    is_curtains[curtain_290]=True
    is_curtain[curtain_290]=True
    is_curtains[curtain_291]=True
    is_curtain[curtain_291]=True
    is_hanger[hanger_292]=True
    is_coatrack[hanger_292]=True
    is_hanger[hanger_293]=True
    is_coatrack[hanger_293]=True
    is_hanger[hanger_294]=True
    is_coatrack[hanger_294]=True
    is_ceilinglamp[ceilinglamp_303]=True
    is_walllamp[walllamp_304]=True
    is_walllamp[walllamp_305]=True
    is_walllamp[walllamp_306]=True
    is_walllamp[walllamp_307]=True
    is_doorjamb[doorjamb_308]=True
    is_doorjamb[doorjamb_309]=True
    is_window[window_310]=True
    is_creamybuns[food_food_1000]=True
    is_cutlets[food_food_1000]=True
    is_salmon[food_food_1000]=True
    is_pear[food_food_1000]=True
    is_chicken[food_food_1000]=True
    is_plum[food_food_1000]=True
    is_orange[food_food_1000]=True
    is_cereal[food_food_1000]=True
    is_banana[food_food_1000]=True
    is_bell_pepper[food_food_1000]=True
    is_apple[food_food_1000]=True
    is_whippedcream[food_food_1000]=True
    is_chinesefood[food_food_1000]=True
    is_food_food[food_food_1000]=True
    is_tomato[food_food_1000]=True
    is_bananas[food_food_1000]=True
    is_chocolatesyrup[food_food_1000]=True
    is_potato[food_food_1000]=True
    is_bellpepper[food_food_1000]=True
    is_crackers[food_food_1000]=True
    is_cucumber[food_food_1000]=True
    is_wooden_spoon[wooden_spoon_2000]=True
    is_creamybuns[food_food_2001]=True
    is_cutlets[food_food_2001]=True
    is_salmon[food_food_2001]=True
    is_pear[food_food_2001]=True
    is_chicken[food_food_2001]=True
    is_plum[food_food_2001]=True
    is_orange[food_food_2001]=True
    is_cereal[food_food_2001]=True
    is_banana[food_food_2001]=True
    is_bell_pepper[food_food_2001]=True
    is_apple[food_food_2001]=True
    is_whippedcream[food_food_2001]=True
    is_chinesefood[food_food_2001]=True
    is_food_food[food_food_2001]=True
    is_tomato[food_food_2001]=True
    is_bananas[food_food_2001]=True
    is_chocolatesyrup[food_food_2001]=True
    is_potato[food_food_2001]=True
    is_bellpepper[food_food_2001]=True
    is_crackers[food_food_2001]=True
    is_cucumber[food_food_2001]=True
    is_brush[brush_2002]=True
    is_chair[chair_2003]=True
    is_lighter[lighter_2004]=True
    is_table_cloth[table_cloth_2005]=True
    is_placemat[table_cloth_2005]=True
    is_piano_bench[piano_bench_2006]=True
    is_food_butter[food_butter_2007]=True
    is_journal[diary_2008]=True
    is_diary[diary_2008]=True
    is_food_onion[food_onion_2009]=True
    is_soap[soap_2010]=True
    is_barsoap[soap_2010]=True
    is_dishwashingliquid[detergent_2011]=True
    is_detergent[detergent_2011]=True
    is_measuring_cup[measuring_cup_2012]=True
    is_oil[oil_2013]=True
    is_condiment_bottle[oil_2013]=True
    is_pen[pencil_2014]=True
    is_pencil[pencil_2014]=True
    is_food_carrot[food_carrot_2015]=True
    is_carrot[food_carrot_2015]=True
    is_wall_phone[phone_2016]=True
    is_phone[phone_2016]=True
    is_cellphone[phone_2016]=True
    is_wall_phone[phone_2017]=True
    is_phone[phone_2017]=True
    is_cellphone[phone_2017]=True
    is_envelope[envelope_2018]=True
    is_hairproduct[shampoo_2019]=True
    is_shampoo[shampoo_2019]=True
    is_lotionbottle[shampoo_2019]=True
    is_pen[pencil_2020]=True
    is_pencil[pencil_2020]=True
    is_creamybuns[food_food_2021]=True
    is_cutlets[food_food_2021]=True
    is_salmon[food_food_2021]=True
    is_pear[food_food_2021]=True
    is_chicken[food_food_2021]=True
    is_plum[food_food_2021]=True
    is_orange[food_food_2021]=True
    is_cereal[food_food_2021]=True
    is_banana[food_food_2021]=True
    is_bell_pepper[food_food_2021]=True
    is_apple[food_food_2021]=True
    is_whippedcream[food_food_2021]=True
    is_chinesefood[food_food_2021]=True
    is_food_food[food_food_2021]=True
    is_tomato[food_food_2021]=True
    is_bananas[food_food_2021]=True
    is_chocolatesyrup[food_food_2021]=True
    is_potato[food_food_2021]=True
    is_bellpepper[food_food_2021]=True
    is_crackers[food_food_2021]=True
    is_cucumber[food_food_2021]=True
    is_stamp[stamp_2022]=True
    is_tea_bag[tea_bag_2023]=True
    is_ice[ice_2024]=True
    is_rag[rag_2025]=True
    is_paper[check_2026]=True
    is_check[check_2026]=True
    is_food_orange[food_orange_2027]=True
    is_instrument_guitar[instrument_guitar_2028]=True
    is_wall_phone[phone_2029]=True
    is_phone[phone_2029]=True
    is_cellphone[phone_2029]=True
    is_cd[cd_2030]=True
    is_scrabble[scrabble_2031]=True
    is_slippers[shoes_2033]=True
    is_shoes[shoes_2033]=True
    is_laser_pointer[laser_pointer_2034]=True
    is_chefknife[knife_2035]=True
    is_cutlery_knife[knife_2035]=True
    is_knife[knife_2035]=True
    is_pants[clothes_pants_2036]=True
    is_clothes_pants[clothes_pants_2036]=True
    is_chefknife[knife_2037]=True
    is_cutlery_knife[knife_2037]=True
    is_knife[knife_2037]=True
    is_box[box_2038]=True
    is_lighter[lighter_2039]=True
    is_pot[pot_2040]=True
    is_condiment_shaker[food_salt_2041]=True
    is_food_salt[food_salt_2041]=True
    is_face_cream[after_shave_2042]=True
    is_facecream[after_shave_2042]=True
    is_after_shave[after_shave_2042]=True
    is_stamp[stamp_2043]=True
    is_shoe_rack[shoe_rack_2044]=True
    is_glue[glue_2045]=True
    is_creamybuns[food_food_2046]=True
    is_cutlets[food_food_2046]=True
    is_salmon[food_food_2046]=True
    is_pear[food_food_2046]=True
    is_chicken[food_food_2046]=True
    is_plum[food_food_2046]=True
    is_orange[food_food_2046]=True
    is_cereal[food_food_2046]=True
    is_banana[food_food_2046]=True
    is_bell_pepper[food_food_2046]=True
    is_apple[food_food_2046]=True
    is_whippedcream[food_food_2046]=True
    is_chinesefood[food_food_2046]=True
    is_food_food[food_food_2046]=True
    is_tomato[food_food_2046]=True
    is_bananas[food_food_2046]=True
    is_chocolatesyrup[food_food_2046]=True
    is_potato[food_food_2046]=True
    is_bellpepper[food_food_2046]=True
    is_crackers[food_food_2046]=True
    is_cucumber[food_food_2046]=True
    is_homework[homework_2047]=True
    is_food_onion[food_onion_2048]=True
    is_wineglass[cup_2049]=True
    is_cup[cup_2049]=True
    is_waterglass[cup_2049]=True
    is_mug[cup_2049]=True
    is_stereo[stereo_2050]=True
    is_radio[stereo_2050]=True
    is_face_cream[after_shave_2051]=True
    is_facecream[after_shave_2051]=True
    is_after_shave[after_shave_2051]=True
    is_rag[rag_2052]=True
    is_coffee_filter[coffee_filter_2053]=True
    is_food_kiwi[food_kiwi_2054]=True
    is_envelope[envelope_2055]=True
    is_sportsball[toy_2056]=True
    is_teddybear[toy_2056]=True
    is_globe[toy_2056]=True
    is_toy[toy_2056]=True
    is_blow_dryer[blow_dryer_2057]=True
    is_paper[check_2058]=True
    is_check[check_2058]=True
    is_toothpaste[tooth_paste_2059]=True
    is_tooth_paste[tooth_paste_2059]=True
    is_book[novel_2060]=True
    is_novel[novel_2060]=True
    is_food_orange[food_orange_2061]=True
    is_piano_bench[piano_bench_2062]=True
    is_face_cream[after_shave_2063]=True
    is_facecream[after_shave_2063]=True
    is_after_shave[after_shave_2063]=True
    is_creamybuns[food_food_2064]=True
    is_cutlets[food_food_2064]=True
    is_salmon[food_food_2064]=True
    is_pear[food_food_2064]=True
    is_chicken[food_food_2064]=True
    is_plum[food_food_2064]=True
    is_orange[food_food_2064]=True
    is_cereal[food_food_2064]=True
    is_banana[food_food_2064]=True
    is_bell_pepper[food_food_2064]=True
    is_apple[food_food_2064]=True
    is_whippedcream[food_food_2064]=True
    is_chinesefood[food_food_2064]=True
    is_food_food[food_food_2064]=True
    is_tomato[food_food_2064]=True
    is_bananas[food_food_2064]=True
    is_chocolatesyrup[food_food_2064]=True
    is_potato[food_food_2064]=True
    is_bellpepper[food_food_2064]=True
    is_crackers[food_food_2064]=True
    is_cucumber[food_food_2064]=True
    is_coffee_filter[coffee_filter_2065]=True
    is_tea[tea_2066]=True
    is_piano_bench[piano_bench_2067]=True
    is_oventray[tray_2068]=True
    is_tray[tray_2068]=True
    is_cat[cat_2069]=True
    is_chessboard[chessboard_2070]=True
    is_paper[check_2071]=True
    is_check[check_2071]=True
    is_food_cheese[food_cheese_2072]=True
    is_creamybuns[food_food_2073]=True
    is_cutlets[food_food_2073]=True
    is_salmon[food_food_2073]=True
    is_pear[food_food_2073]=True
    is_chicken[food_food_2073]=True
    is_plum[food_food_2073]=True
    is_orange[food_food_2073]=True
    is_cereal[food_food_2073]=True
    is_banana[food_food_2073]=True
    is_bell_pepper[food_food_2073]=True
    is_apple[food_food_2073]=True
    is_whippedcream[food_food_2073]=True
    is_chinesefood[food_food_2073]=True
    is_food_food[food_food_2073]=True
    is_tomato[food_food_2073]=True
    is_bananas[food_food_2073]=True
    is_chocolatesyrup[food_food_2073]=True
    is_potato[food_food_2073]=True
    is_bellpepper[food_food_2073]=True
    is_crackers[food_food_2073]=True
    is_cucumber[food_food_2073]=True
    is_creamybuns[food_food_2074]=True
    is_cutlets[food_food_2074]=True
    is_salmon[food_food_2074]=True
    is_pear[food_food_2074]=True
    is_chicken[food_food_2074]=True
    is_plum[food_food_2074]=True
    is_orange[food_food_2074]=True
    is_cereal[food_food_2074]=True
    is_banana[food_food_2074]=True
    is_bell_pepper[food_food_2074]=True
    is_apple[food_food_2074]=True
    is_whippedcream[food_food_2074]=True
    is_chinesefood[food_food_2074]=True
    is_food_food[food_food_2074]=True
    is_tomato[food_food_2074]=True
    is_bananas[food_food_2074]=True
    is_chocolatesyrup[food_food_2074]=True
    is_potato[food_food_2074]=True
    is_bellpepper[food_food_2074]=True
    is_crackers[food_food_2074]=True
    is_cucumber[food_food_2074]=True
    is_paper[check_2075]=True
    is_check[check_2075]=True
    is_toiletpaper[toilet_paper_2076]=True
    is_toilet_paper[toilet_paper_2076]=True
    is_food_peanut_butter[food_peanut_butter_2077]=True
    #categories_end

    #states
    is_on[walllamp_34]=True
    is_on[ceilinglamp_35]=True
    is_on[walllamp_36]=True
    is_on[fridge_126]=True
    is_on[toaster_132]=True
    is_on[ceilinglamp_137]=True
    is_on[ceilinglamp_138]=True
    is_on[walllamp_139]=True
    is_on[walllamp_140]=True
    is_on[walllamp_141]=True
    is_on[ceilinglamp_237]=True
    is_on[tablelamp_238]=True
    is_on[tablelamp_239]=True
    is_on[ceilinglamp_303]=True
    is_on[walllamp_304]=True
    is_on[walllamp_305]=True
    is_on[walllamp_306]=True
    is_on[walllamp_307]=True
    is_on[lighter_2004]=True
    is_on[laser_pointer_2034]=True
    is_on[lighter_2039]=True
    is_off[iron_2161]=True
    is_off[washing_machine_2079]=True
    is_off[remote_control_2124]=True
    is_off[cd_player_2129]=True
    is_off[dvd_player_2130]=True
    is_off[stove_2135]=True
    is_off[vacuum_cleaner_2139]=True
    is_off[phone_2147]=True
    is_off[toilet_15]=True
    is_off[faucet_20]=True
    is_off[light_39]=True
    is_off[phone_71]=True
    is_off[light_73]=True
    is_off[faucet_121]=True
    is_off[oven_127]=True
    is_off[dishwasher_129]=True
    is_off[coffe_maker_130]=True
    is_off[microwave_135]=True
    is_off[computer_209]=True
    is_off[light_212]=True
    is_off[computer_276]=True
    is_off[television_281]=True
    is_off[light_283]=True
    is_off[phone_2017]=True
    is_off[instrument_guitar_2028]=True
    is_off[blow_dryer_2057]=True
    open[basket_for_clothes_2078]=True
    open[doorjamb_37]=True
    open[door_38]=True
    open[door_61]=True
    open[door_62]=True
    open[pot_78]=True
    open[trashcan_99]=True
    open[cupboard_117]=True
    open[kitchen_counter_119]=True
    open[doorjamb_190]=True
    open[nightstand_192]=True
    open[curtain_206]=True
    open[bookshelf_275]=True
    open[curtain_289]=True
    open[curtain_290]=True
    open[doorjamb_308]=True
    open[doorjamb_309]=True
    open[envelope_2018]=True
    open[shampoo_2019]=True
    open[box_2038]=True
    open[after_shave_2063]=True
    closed[washing_machine_2079]=True
    closed[cd_player_2129]=True
    closed[dvd_player_2130]=True
    closed[stove_2135]=True
    closed[book_2136]=True
    closed[book_2137]=True
    closed[pot_2138]=True
    closed[window_2156]=True
    closed[toilet_15]=True
    closed[bathroom_cabinet_17]=True
    closed[bathroom_counter_18]=True
    closed[curtain_22]=True
    closed[light_39]=True
    closed[light_73]=True
    closed[cupboard_118]=True
    closed[kitchen_counter_122]=True
    closed[kitchen_counter_123]=True
    closed[bookshelf_124]=True
    closed[fridge_126]=True
    closed[oven_127]=True
    closed[dishwasher_129]=True
    closed[coffe_maker_130]=True
    closed[microwave_135]=True
    closed[window_191]=True
    closed[nightstand_195]=True
    closed[bookshelf_196]=True
    closed[filing_cabinet_200]=True
    closed[curtain_204]=True
    closed[curtain_205]=True
    closed[light_212]=True
    closed[desk_272]=True
    closed[dresser_274]=True
    closed[light_283]=True
    closed[curtain_291]=True
    closed[window_310]=True
    closed[diary_2008]=True
    closed[pot_2040]=True
    closed[after_shave_2042]=True
    closed[stereo_2050]=True
    closed[after_shave_2051]=True
    closed[envelope_2055]=True
    closed[tooth_paste_2059]=True
    closed[novel_2060]=True
    dirty[clothes_pants_2157]=True
    dirty[clothes_shirt_2158]=True
    dirty[clothes_socks_2159]=True
    dirty[clothes_skirt_2160]=True
    dirty[food_vegetable_2113]=True
    dirty[clothes_dress_2116]=True
    dirty[clothes_jacket_2119]=True
    dirty[clothes_scarf_2120]=True
    dirty[clothes_underwear_2121]=True
    dirty[bowl_2140]=True
    dirty[bowl_2141]=True
    dirty[bowl_2142]=True
    dirty[plate_2152]=True
    dirty[window_2156]=True
    dirty[wall_2]=True
    dirty[wall_5]=True
    dirty[floor_10]=True
    dirty[floor_12]=True
    dirty[floor_13]=True
    dirty[floor_14]=True
    dirty[sink_19]=True
    dirty[floor_43]=True
    dirty[floor_47]=True
    dirty[floor_49]=True
    dirty[floor_51]=True
    dirty[ceiling_53]=True
    dirty[ceiling_55]=True
    dirty[ceiling_56]=True
    dirty[ceiling_58]=True
    dirty[ceiling_59]=True
    dirty[ceiling_60]=True
    dirty[wall_63]=True
    dirty[wall_64]=True
    dirty[wall_66]=True
    dirty[wall_68]=True
    dirty[wall_70]=True
    dirty[pillow_104]=True
    dirty[pillow_105]=True
    dirty[table_114]=True
    dirty[sink_120]=True
    dirty[kitchen_counter_122]=True
    dirty[tray_128]=True
    dirty[microwave_135]=True
    dirty[floor_165]=True
    dirty[floor_168]=True
    dirty[floor_169]=True
    dirty[floor_170]=True
    dirty[floor_171]=True
    dirty[floor_172]=True
    dirty[wall_173]=True
    dirty[wall_178]=True
    dirty[wall_179]=True
    dirty[wall_180]=True
    dirty[ceiling_181]=True
    dirty[ceiling_183]=True
    dirty[ceiling_184]=True
    dirty[ceiling_186]=True
    dirty[window_191]=True
    dirty[bookshelf_196]=True
    dirty[table_199]=True
    dirty[filing_cabinet_200]=True
    dirty[curtain_204]=True
    dirty[pillow_207]=True
    dirty[wall_242]=True
    dirty[wall_243]=True
    dirty[wall_244]=True
    dirty[wall_245]=True
    dirty[wall_248]=True
    dirty[wall_249]=True
    dirty[ceiling_251]=True
    dirty[ceiling_252]=True
    dirty[ceiling_254]=True
    dirty[ceiling_257]=True
    dirty[ceiling_258]=True
    dirty[floor_259]=True
    dirty[floor_260]=True
    dirty[floor_262]=True
    dirty[floor_264]=True
    dirty[floor_265]=True
    dirty[mousepad_279]=True
    dirty[curtain_291]=True
    dirty[window_310]=True
    dirty[wooden_spoon_2000]=True
    dirty[food_food_2001]=True
    dirty[food_carrot_2015]=True
    dirty[food_food_2021]=True
    dirty[food_orange_2027]=True
    dirty[cd_2030]=True
    dirty[food_food_2046]=True
    dirty[cup_2049]=True
    dirty[coffee_filter_2053]=True
    dirty[piano_bench_2062]=True
    dirty[food_food_2064]=True
    dirty[food_food_2073]=True
    clean[iron_2161]=True
    clean[washing_machine_2079]=True
    clean[food_steak_2080]=True
    clean[food_apple_2081]=True
    clean[food_bacon_2082]=True
    clean[food_banana_2083]=True
    clean[food_bread_2084]=True
    clean[food_cake_2085]=True
    clean[food_carrot_2086]=True
    clean[food_cereal_2087]=True
    clean[food_cheese_2088]=True
    clean[food_chicken_2089]=True
    clean[food_dessert_2090]=True
    clean[food_donut_2091]=True
    clean[food_egg_2092]=True
    clean[food_fish_2093]=True
    clean[food_food_2094]=True
    clean[food_fruit_2095]=True
    clean[food_hamburger_2096]=True
    clean[food_ice_cream_2097]=True
    clean[food_jam_2098]=True
    clean[food_kiwi_2099]=True
    clean[food_lemon_2100]=True
    clean[food_noodles_2101]=True
    clean[food_oatmeal_2102]=True
    clean[food_orange_2103]=True
    clean[food_onion_2104]=True
    clean[food_peanut_butter_2105]=True
    clean[food_pizza_2106]=True
    clean[food_potato_2107]=True
    clean[food_rice_2108]=True
    clean[food_salt_2109]=True
    clean[food_snack_2110]=True
    clean[food_sugar_2111]=True
    clean[food_turkey_2112]=True
    clean[dry_pasta_2114]=True
    clean[clothes_hat_2117]=True
    clean[clothes_gloves_2118]=True
    clean[knife_2122]=True
    clean[cutting_board_2123]=True
    clean[soap_2125]=True
    clean[soap_2126]=True
    clean[towel_2128]=True
    clean[vacuum_cleaner_2139]=True
    clean[phone_2147]=True
    clean[fork_2150]=True
    clean[fork_2151]=True
    clean[fryingpan_2154]=True
    clean[detergent_2155]=True
    clean[bathroom_1]=True
    clean[wall_3]=True
    clean[wall_4]=True
    clean[ceiling_6]=True
    clean[ceiling_7]=True
    clean[ceiling_8]=True
    clean[ceiling_9]=True
    clean[floor_11]=True
    clean[toilet_15]=True
    clean[shower_16]=True
    clean[bathroom_cabinet_17]=True
    clean[bathroom_counter_18]=True
    clean[faucet_20]=True
    clean[shower_21]=True
    clean[curtain_22]=True
    clean[mat_32]=True
    clean[drawing_33]=True
    clean[walllamp_34]=True
    clean[ceilinglamp_35]=True
    clean[walllamp_36]=True
    clean[doorjamb_37]=True
    clean[door_38]=True
    clean[light_39]=True
    clean[dining_room_41]=True
    clean[floor_42]=True
    clean[floor_44]=True
    clean[floor_45]=True
    clean[floor_46]=True
    clean[floor_48]=True
    clean[floor_50]=True
    clean[ceiling_52]=True
    clean[ceiling_54]=True
    clean[ceiling_57]=True
    clean[door_61]=True
    clean[door_62]=True
    clean[wall_65]=True
    clean[wall_67]=True
    clean[wall_69]=True
    clean[phone_71]=True
    clean[powersocket_72]=True
    clean[light_73]=True
    clean[knifeblock_76]=True
    clean[pot_78]=True
    clean[trashcan_99]=True
    clean[mat_102]=True
    clean[pillow_103]=True
    clean[pillow_106]=True
    clean[pillow_107]=True
    clean[pillow_108]=True
    clean[drawing_110]=True
    clean[drawing_111]=True
    clean[bench_113]=True
    clean[bench_115]=True
    clean[tvstand_116]=True
    clean[cupboard_117]=True
    clean[cupboard_118]=True
    clean[kitchen_counter_119]=True
    clean[faucet_121]=True
    clean[kitchen_counter_123]=True
    clean[bookshelf_124]=True
    clean[stovefan_125]=True
    clean[fridge_126]=True
    clean[oven_127]=True
    clean[dishwasher_129]=True
    clean[coffe_maker_130]=True
    clean[toaster_132]=True
    clean[ceilinglamp_137]=True
    clean[ceilinglamp_138]=True
    clean[walllamp_139]=True
    clean[walllamp_140]=True
    clean[walllamp_141]=True
    clean[bedroom_162]=True
    clean[floor_163]=True
    clean[floor_164]=True
    clean[floor_166]=True
    clean[floor_167]=True
    clean[wall_174]=True
    clean[wall_175]=True
    clean[wall_176]=True
    clean[wall_177]=True
    clean[ceiling_182]=True
    clean[ceiling_185]=True
    clean[ceiling_187]=True
    clean[ceiling_188]=True
    clean[ceiling_189]=True
    clean[doorjamb_190]=True
    clean[nightstand_192]=True
    clean[desk_193]=True
    clean[chair_194]=True
    clean[nightstand_195]=True
    clean[bed_197]=True
    clean[couch_198]=True
    clean[drawing_201]=True
    clean[drawing_202]=True
    clean[mat_203]=True
    clean[curtain_205]=True
    clean[curtain_206]=True
    clean[pillow_208]=True
    clean[computer_209]=True
    clean[cpuscreen_210]=True
    clean[keyboard_211]=True
    clean[light_212]=True
    clean[mouse_213]=True
    clean[mousepad_214]=True
    clean[photoframe_219]=True
    clean[ceilinglamp_237]=True
    clean[tablelamp_238]=True
    clean[tablelamp_239]=True
    clean[home_office_241]=True
    clean[wall_246]=True
    clean[wall_247]=True
    clean[ceiling_250]=True
    clean[ceiling_253]=True
    clean[ceiling_255]=True
    clean[ceiling_256]=True
    clean[floor_261]=True
    clean[floor_263]=True
    clean[floor_266]=True
    clean[floor_267]=True
    clean[floor_268]=True
    clean[couch_269]=True
    clean[table_270]=True
    clean[chair_271]=True
    clean[desk_272]=True
    clean[tvstand_273]=True
    clean[dresser_274]=True
    clean[bookshelf_275]=True
    clean[computer_276]=True
    clean[cpuscreen_277]=True
    clean[keyboard_278]=True
    clean[mouse_280]=True
    clean[television_281]=True
    clean[powersocket_282]=True
    clean[light_283]=True
    clean[mat_284]=True
    clean[orchid_285]=True
    clean[pillow_286]=True
    clean[pillow_287]=True
    clean[drawing_288]=True
    clean[curtain_289]=True
    clean[curtain_290]=True
    clean[hanger_292]=True
    clean[hanger_293]=True
    clean[hanger_294]=True
    clean[ceilinglamp_303]=True
    clean[walllamp_304]=True
    clean[walllamp_305]=True
    clean[walllamp_306]=True
    clean[walllamp_307]=True
    clean[doorjamb_308]=True
    clean[doorjamb_309]=True
    clean[food_food_1000]=True
    clean[brush_2002]=True
    clean[chair_2003]=True
    clean[lighter_2004]=True
    clean[table_cloth_2005]=True
    clean[piano_bench_2006]=True
    clean[food_butter_2007]=True
    clean[diary_2008]=True
    clean[food_onion_2009]=True
    clean[soap_2010]=True
    clean[detergent_2011]=True
    clean[measuring_cup_2012]=True
    clean[oil_2013]=True
    clean[pencil_2014]=True
    clean[phone_2016]=True
    clean[phone_2017]=True
    clean[envelope_2018]=True
    clean[shampoo_2019]=True
    clean[pencil_2020]=True
    clean[stamp_2022]=True
    clean[tea_bag_2023]=True
    clean[ice_2024]=True
    clean[rag_2025]=True
    clean[check_2026]=True
    clean[instrument_guitar_2028]=True
    clean[phone_2029]=True
    clean[scrabble_2031]=True
    clean[shoes_2033]=True
    clean[laser_pointer_2034]=True
    clean[knife_2035]=True
    clean[clothes_pants_2036]=True
    clean[knife_2037]=True
    clean[box_2038]=True
    clean[lighter_2039]=True
    clean[pot_2040]=True
    clean[food_salt_2041]=True
    clean[after_shave_2042]=True
    clean[stamp_2043]=True
    clean[shoe_rack_2044]=True
    clean[glue_2045]=True
    clean[homework_2047]=True
    clean[food_onion_2048]=True
    clean[stereo_2050]=True
    clean[after_shave_2051]=True
    clean[rag_2052]=True
    clean[food_kiwi_2054]=True
    clean[envelope_2055]=True
    clean[toy_2056]=True
    clean[blow_dryer_2057]=True
    clean[check_2058]=True
    clean[tooth_paste_2059]=True
    clean[novel_2060]=True
    clean[food_orange_2061]=True
    clean[after_shave_2063]=True
    clean[coffee_filter_2065]=True
    clean[tea_2066]=True
    clean[piano_bench_2067]=True
    clean[tray_2068]=True
    clean[cat_2069]=True
    clean[chessboard_2070]=True
    clean[check_2071]=True
    clean[food_cheese_2072]=True
    clean[food_food_2074]=True
    clean[check_2075]=True
    clean[toilet_paper_2076]=True
    clean[food_peanut_butter_2077]=True
    plugged[light_39]=True
    plugged[phone_71]=True
    plugged[light_73]=True
    plugged[fridge_126]=True
    plugged[oven_127]=True
    plugged[dishwasher_129]=True
    plugged[coffe_maker_130]=True
    plugged[toaster_132]=True
    plugged[microwave_135]=True
    plugged[computer_209]=True
    plugged[keyboard_211]=True
    plugged[light_212]=True
    plugged[computer_276]=True
    plugged[keyboard_278]=True
    plugged[television_281]=True
    plugged[light_283]=True
    plugged[phone_2017]=True
    plugged[blow_dryer_2057]=True
    unplugged[iron_2161]=True
    unplugged[washing_machine_2079]=True
    unplugged[cd_player_2129]=True
    unplugged[dvd_player_2130]=True
    unplugged[vacuum_cleaner_2139]=True
    unplugged[mouse_213]=True
    unplugged[mouse_280]=True
    unplugged[phone_2016]=True
    unplugged[phone_2029]=True
    unplugged[stereo_2050]=True
    is_room[bathroom_1]=True
    is_room[dining_room_41]=True
    is_room[bedroom_162]=True
    is_room[home_office_241]=True
    #states_end

    #char_states
    standing[char]=True
    sitting[char]=False
    lying[char]=False
    sleeping[char]=False
    has_a_free_hand[char]=True
    #char_states_end

    #char
    inside_char[char,dining_room_41]=True
    #char_end

    #properties
    surfaces[cutting_board_2123]=True
    surfaces[cd_player_2129]=True
    surfaces[dvd_player_2130]=True
    surfaces[stove_2135]=True
    surfaces[ironing_board_2144]=True
    surfaces[plate_2152]=True
    surfaces[floor_10]=True
    surfaces[floor_11]=True
    surfaces[floor_12]=True
    surfaces[floor_13]=True
    surfaces[floor_14]=True
    surfaces[bathroom_cabinet_17]=True
    surfaces[bathroom_counter_18]=True
    surfaces[mat_32]=True
    surfaces[floor_42]=True
    surfaces[floor_43]=True
    surfaces[floor_44]=True
    surfaces[floor_45]=True
    surfaces[floor_46]=True
    surfaces[floor_47]=True
    surfaces[floor_48]=True
    surfaces[floor_49]=True
    surfaces[floor_50]=True
    surfaces[floor_51]=True
    surfaces[mat_102]=True
    surfaces[bench_113]=True
    surfaces[table_114]=True
    surfaces[bench_115]=True
    surfaces[tvstand_116]=True
    surfaces[kitchen_counter_119]=True
    surfaces[kitchen_counter_122]=True
    surfaces[kitchen_counter_123]=True
    surfaces[bookshelf_124]=True
    surfaces[tray_128]=True
    surfaces[floor_163]=True
    surfaces[floor_164]=True
    surfaces[floor_165]=True
    surfaces[floor_166]=True
    surfaces[floor_167]=True
    surfaces[floor_168]=True
    surfaces[floor_169]=True
    surfaces[floor_170]=True
    surfaces[floor_171]=True
    surfaces[floor_172]=True
    surfaces[nightstand_192]=True
    surfaces[desk_193]=True
    surfaces[chair_194]=True
    surfaces[nightstand_195]=True
    surfaces[bookshelf_196]=True
    surfaces[bed_197]=True
    surfaces[couch_198]=True
    surfaces[table_199]=True
    surfaces[filing_cabinet_200]=True
    surfaces[mat_203]=True
    surfaces[mousepad_214]=True
    surfaces[floor_259]=True
    surfaces[floor_260]=True
    surfaces[floor_261]=True
    surfaces[floor_262]=True
    surfaces[floor_263]=True
    surfaces[floor_264]=True
    surfaces[floor_265]=True
    surfaces[floor_266]=True
    surfaces[floor_267]=True
    surfaces[floor_268]=True
    surfaces[couch_269]=True
    surfaces[table_270]=True
    surfaces[chair_271]=True
    surfaces[desk_272]=True
    surfaces[tvstand_273]=True
    surfaces[bookshelf_275]=True
    surfaces[mousepad_279]=True
    surfaces[mat_284]=True
    surfaces[chair_2003]=True
    surfaces[table_cloth_2005]=True
    surfaces[piano_bench_2006]=True
    surfaces[shoe_rack_2044]=True
    surfaces[stereo_2050]=True
    surfaces[piano_bench_2062]=True
    surfaces[piano_bench_2067]=True
    surfaces[tray_2068]=True
    surfaces[chessboard_2070]=True
    grabbable[clothes_pants_2157]=True
    grabbable[clothes_shirt_2158]=True
    grabbable[clothes_socks_2159]=True
    grabbable[clothes_skirt_2160]=True
    grabbable[iron_2161]=True
    grabbable[basket_for_clothes_2078]=True
    grabbable[food_steak_2080]=True
    grabbable[food_apple_2081]=True
    grabbable[food_bacon_2082]=True
    grabbable[food_banana_2083]=True
    grabbable[food_bread_2084]=True
    grabbable[food_cake_2085]=True
    grabbable[food_carrot_2086]=True
    grabbable[food_cereal_2087]=True
    grabbable[food_cheese_2088]=True
    grabbable[food_chicken_2089]=True
    grabbable[food_dessert_2090]=True
    grabbable[food_donut_2091]=True
    grabbable[food_egg_2092]=True
    grabbable[food_fish_2093]=True
    grabbable[food_food_2094]=True
    grabbable[food_fruit_2095]=True
    grabbable[food_hamburger_2096]=True
    grabbable[food_ice_cream_2097]=True
    grabbable[food_jam_2098]=True
    grabbable[food_kiwi_2099]=True
    grabbable[food_lemon_2100]=True
    grabbable[food_noodles_2101]=True
    grabbable[food_oatmeal_2102]=True
    grabbable[food_orange_2103]=True
    grabbable[food_onion_2104]=True
    grabbable[food_peanut_butter_2105]=True
    grabbable[food_pizza_2106]=True
    grabbable[food_potato_2107]=True
    grabbable[food_rice_2108]=True
    grabbable[food_salt_2109]=True
    grabbable[food_snack_2110]=True
    grabbable[food_sugar_2111]=True
    grabbable[food_turkey_2112]=True
    grabbable[food_vegetable_2113]=True
    grabbable[dry_pasta_2114]=True
    grabbable[milk_2115]=True
    grabbable[clothes_dress_2116]=True
    grabbable[clothes_hat_2117]=True
    grabbable[clothes_gloves_2118]=True
    grabbable[clothes_jacket_2119]=True
    grabbable[clothes_scarf_2120]=True
    grabbable[clothes_underwear_2121]=True
    grabbable[knife_2122]=True
    grabbable[cutting_board_2123]=True
    grabbable[remote_control_2124]=True
    grabbable[soap_2125]=True
    grabbable[soap_2126]=True
    grabbable[towel_2128]=True
    grabbable[cd_player_2129]=True
    grabbable[dvd_player_2130]=True
    grabbable[headset_2131]=True
    grabbable[cup_2132]=True
    grabbable[cup_2133]=True
    grabbable[cup_2134]=True
    grabbable[book_2136]=True
    grabbable[book_2137]=True
    grabbable[pot_2138]=True
    grabbable[vacuum_cleaner_2139]=True
    grabbable[bowl_2140]=True
    grabbable[bowl_2141]=True
    grabbable[bowl_2142]=True
    grabbable[cleaning_solution_2143]=True
    grabbable[cd_2145]=True
    grabbable[headset_2146]=True
    grabbable[phone_2147]=True
    grabbable[sauce_2148]=True
    grabbable[oil_2149]=True
    grabbable[fork_2150]=True
    grabbable[fork_2151]=True
    grabbable[plate_2152]=True
    grabbable[spectacles_2153]=True
    grabbable[fryingpan_2154]=True
    grabbable[detergent_2155]=True
    grabbable[mat_32]=True
    grabbable[drawing_33]=True
    grabbable[phone_71]=True
    grabbable[pot_78]=True
    grabbable[mat_102]=True
    grabbable[pillow_103]=True
    grabbable[pillow_104]=True
    grabbable[pillow_105]=True
    grabbable[pillow_106]=True
    grabbable[pillow_107]=True
    grabbable[pillow_108]=True
    grabbable[drawing_110]=True
    grabbable[drawing_111]=True
    grabbable[tray_128]=True
    grabbable[chair_194]=True
    grabbable[drawing_201]=True
    grabbable[drawing_202]=True
    grabbable[mat_203]=True
    grabbable[pillow_207]=True
    grabbable[pillow_208]=True
    grabbable[keyboard_211]=True
    grabbable[mouse_213]=True
    grabbable[chair_271]=True
    grabbable[keyboard_278]=True
    grabbable[mouse_280]=True
    grabbable[mat_284]=True
    grabbable[pillow_286]=True
    grabbable[pillow_287]=True
    grabbable[drawing_288]=True
    grabbable[hanger_292]=True
    grabbable[hanger_293]=True
    grabbable[hanger_294]=True
    grabbable[food_food_1000]=True
    grabbable[wooden_spoon_2000]=True
    grabbable[food_food_2001]=True
    grabbable[brush_2002]=True
    grabbable[chair_2003]=True
    grabbable[lighter_2004]=True
    grabbable[table_cloth_2005]=True
    grabbable[piano_bench_2006]=True
    grabbable[food_butter_2007]=True
    grabbable[diary_2008]=True
    grabbable[food_onion_2009]=True
    grabbable[soap_2010]=True
    grabbable[detergent_2011]=True
    grabbable[measuring_cup_2012]=True
    grabbable[oil_2013]=True
    grabbable[pencil_2014]=True
    grabbable[food_carrot_2015]=True
    grabbable[phone_2016]=True
    grabbable[phone_2017]=True
    grabbable[envelope_2018]=True
    grabbable[shampoo_2019]=True
    grabbable[pencil_2020]=True
    grabbable[food_food_2021]=True
    grabbable[stamp_2022]=True
    grabbable[tea_bag_2023]=True
    grabbable[ice_2024]=True
    grabbable[rag_2025]=True
    grabbable[check_2026]=True
    grabbable[food_orange_2027]=True
    grabbable[instrument_guitar_2028]=True
    grabbable[phone_2029]=True
    grabbable[cd_2030]=True
    grabbable[scrabble_2031]=True
    grabbable[shoes_2033]=True
    grabbable[laser_pointer_2034]=True
    grabbable[knife_2035]=True
    grabbable[clothes_pants_2036]=True
    grabbable[knife_2037]=True
    grabbable[box_2038]=True
    grabbable[lighter_2039]=True
    grabbable[pot_2040]=True
    grabbable[food_salt_2041]=True
    grabbable[after_shave_2042]=True
    grabbable[stamp_2043]=True
    grabbable[shoe_rack_2044]=True
    grabbable[glue_2045]=True
    grabbable[food_food_2046]=True
    grabbable[homework_2047]=True
    grabbable[food_onion_2048]=True
    grabbable[cup_2049]=True
    grabbable[stereo_2050]=True
    grabbable[after_shave_2051]=True
    grabbable[rag_2052]=True
    grabbable[coffee_filter_2053]=True
    grabbable[food_kiwi_2054]=True
    grabbable[envelope_2055]=True
    grabbable[toy_2056]=True
    grabbable[blow_dryer_2057]=True
    grabbable[check_2058]=True
    grabbable[tooth_paste_2059]=True
    grabbable[novel_2060]=True
    grabbable[food_orange_2061]=True
    grabbable[piano_bench_2062]=True
    grabbable[after_shave_2063]=True
    grabbable[food_food_2064]=True
    grabbable[coffee_filter_2065]=True
    grabbable[tea_2066]=True
    grabbable[piano_bench_2067]=True
    grabbable[tray_2068]=True
    grabbable[cat_2069]=True
    grabbable[chessboard_2070]=True
    grabbable[check_2071]=True
    grabbable[food_cheese_2072]=True
    grabbable[food_food_2073]=True
    grabbable[food_food_2074]=True
    grabbable[check_2075]=True
    grabbable[toilet_paper_2076]=True
    grabbable[food_peanut_butter_2077]=True
    sittable[toilet_15]=True
    sittable[mat_32]=True
    sittable[mat_102]=True
    sittable[bench_113]=True
    sittable[bench_115]=True
    sittable[chair_194]=True
    sittable[bed_197]=True
    sittable[couch_198]=True
    sittable[mat_203]=True
    sittable[couch_269]=True
    sittable[chair_271]=True
    sittable[mat_284]=True
    sittable[chair_2003]=True
    sittable[piano_bench_2006]=True
    sittable[piano_bench_2062]=True
    sittable[piano_bench_2067]=True
    lieable[mat_32]=True
    lieable[mat_102]=True
    lieable[bench_113]=True
    lieable[bench_115]=True
    lieable[bed_197]=True
    lieable[couch_198]=True
    lieable[mat_203]=True
    lieable[couch_269]=True
    lieable[mat_284]=True
    hangable[clothes_pants_2157]=True
    hangable[clothes_shirt_2158]=True
    hangable[clothes_socks_2159]=True
    hangable[clothes_skirt_2160]=True
    hangable[clothes_dress_2116]=True
    hangable[clothes_hat_2117]=True
    hangable[clothes_gloves_2118]=True
    hangable[clothes_jacket_2119]=True
    hangable[clothes_scarf_2120]=True
    hangable[clothes_underwear_2121]=True
    hangable[hanger_292]=True
    hangable[hanger_293]=True
    hangable[hanger_294]=True
    hangable[clothes_pants_2036]=True
    hangable[toilet_paper_2076]=True
    drinkable[milk_2115]=True
    drinkable[oil_2149]=True
    drinkable[oil_2013]=True
    drinkable[tea_2066]=True
    eatable[food_steak_2080]=True
    eatable[food_apple_2081]=True
    eatable[food_bacon_2082]=True
    eatable[food_banana_2083]=True
    eatable[food_bread_2084]=True
    eatable[food_cake_2085]=True
    eatable[food_carrot_2086]=True
    eatable[food_cereal_2087]=True
    eatable[food_cheese_2088]=True
    eatable[food_chicken_2089]=True
    eatable[food_dessert_2090]=True
    eatable[food_egg_2092]=True
    eatable[food_fish_2093]=True
    eatable[food_food_2094]=True
    eatable[food_fruit_2095]=True
    eatable[food_hamburger_2096]=True
    eatable[food_jam_2098]=True
    eatable[food_kiwi_2099]=True
    eatable[food_lemon_2100]=True
    eatable[food_noodles_2101]=True
    eatable[food_oatmeal_2102]=True
    eatable[food_orange_2103]=True
    eatable[food_onion_2104]=True
    eatable[food_peanut_butter_2105]=True
    eatable[food_pizza_2106]=True
    eatable[food_potato_2107]=True
    eatable[food_rice_2108]=True
    eatable[food_salt_2109]=True
    eatable[food_snack_2110]=True
    eatable[food_sugar_2111]=True
    eatable[food_turkey_2112]=True
    eatable[food_vegetable_2113]=True
    eatable[food_food_1000]=True
    eatable[food_food_2001]=True
    eatable[food_onion_2009]=True
    eatable[food_carrot_2015]=True
    eatable[food_food_2021]=True
    eatable[food_orange_2027]=True
    eatable[food_salt_2041]=True
    eatable[food_food_2046]=True
    eatable[food_onion_2048]=True
    eatable[food_kiwi_2054]=True
    eatable[food_orange_2061]=True
    eatable[food_food_2064]=True
    eatable[food_cheese_2072]=True
    eatable[food_food_2073]=True
    eatable[food_food_2074]=True
    eatable[food_peanut_butter_2077]=True
    recipient[washing_machine_2079]=True
    recipient[cup_2132]=True
    recipient[cup_2133]=True
    recipient[cup_2134]=True
    recipient[pot_2138]=True
    recipient[bowl_2140]=True
    recipient[bowl_2141]=True
    recipient[bowl_2142]=True
    recipient[plate_2152]=True
    recipient[fryingpan_2154]=True
    recipient[sink_19]=True
    recipient[pot_78]=True
    recipient[sink_120]=True
    recipient[coffe_maker_130]=True
    recipient[measuring_cup_2012]=True
    recipient[rag_2025]=True
    recipient[box_2038]=True
    recipient[pot_2040]=True
    recipient[cup_2049]=True
    recipient[rag_2052]=True
    cuttable[food_steak_2080]=True
    cuttable[food_apple_2081]=True
    cuttable[food_bacon_2082]=True
    cuttable[food_banana_2083]=True
    cuttable[food_bread_2084]=True
    cuttable[food_cake_2085]=True
    cuttable[food_carrot_2086]=True
    cuttable[food_cheese_2088]=True
    cuttable[food_chicken_2089]=True
    cuttable[food_dessert_2090]=True
    cuttable[food_egg_2092]=True
    cuttable[food_fish_2093]=True
    cuttable[food_food_2094]=True
    cuttable[food_fruit_2095]=True
    cuttable[food_hamburger_2096]=True
    cuttable[food_kiwi_2099]=True
    cuttable[food_lemon_2100]=True
    cuttable[food_orange_2103]=True
    cuttable[food_onion_2104]=True
    cuttable[food_pizza_2106]=True
    cuttable[food_potato_2107]=True
    cuttable[food_turkey_2112]=True
    cuttable[food_vegetable_2113]=True
    cuttable[book_2136]=True
    cuttable[book_2137]=True
    cuttable[drawing_33]=True
    cuttable[drawing_110]=True
    cuttable[drawing_111]=True
    cuttable[drawing_201]=True
    cuttable[drawing_202]=True
    cuttable[drawing_288]=True
    cuttable[food_food_1000]=True
    cuttable[food_food_2001]=True
    cuttable[food_onion_2009]=True
    cuttable[food_carrot_2015]=True
    cuttable[envelope_2018]=True
    cuttable[food_food_2021]=True
    cuttable[food_orange_2027]=True
    cuttable[food_food_2046]=True
    cuttable[food_onion_2048]=True
    cuttable[food_kiwi_2054]=True
    cuttable[envelope_2055]=True
    cuttable[novel_2060]=True
    cuttable[food_orange_2061]=True
    cuttable[food_food_2064]=True
    cuttable[food_cheese_2072]=True
    cuttable[food_food_2073]=True
    cuttable[food_food_2074]=True
    cuttable[toilet_paper_2076]=True
    pourable[food_cereal_2087]=True
    pourable[food_rice_2108]=True
    pourable[food_salt_2109]=True
    pourable[food_sugar_2111]=True
    pourable[milk_2115]=True
    pourable[cup_2132]=True
    pourable[cup_2133]=True
    pourable[cup_2134]=True
    pourable[cleaning_solution_2143]=True
    pourable[sauce_2148]=True
    pourable[oil_2149]=True
    pourable[detergent_2155]=True
    pourable[detergent_2011]=True
    pourable[measuring_cup_2012]=True
    pourable[oil_2013]=True
    pourable[shampoo_2019]=True
    pourable[food_salt_2041]=True
    pourable[after_shave_2042]=True
    pourable[cup_2049]=True
    pourable[after_shave_2051]=True
    pourable[tooth_paste_2059]=True
    pourable[after_shave_2063]=True
    pourable[tea_2066]=True
    can_open[basket_for_clothes_2078]=True
    can_open[washing_machine_2079]=True
    can_open[food_cereal_2087]=True
    can_open[food_jam_2098]=True
    can_open[milk_2115]=True
    can_open[cd_player_2129]=True
    can_open[dvd_player_2130]=True
    can_open[stove_2135]=True
    can_open[book_2136]=True
    can_open[book_2137]=True
    can_open[pot_2138]=True
    can_open[window_2156]=True
    can_open[toilet_15]=True
    can_open[bathroom_cabinet_17]=True
    can_open[curtain_22]=True
    can_open[door_38]=True
    can_open[door_61]=True
    can_open[door_62]=True
    can_open[pot_78]=True
    can_open[trashcan_99]=True
    can_open[cupboard_117]=True
    can_open[cupboard_118]=True
    can_open[bookshelf_124]=True
    can_open[fridge_126]=True
    can_open[oven_127]=True
    can_open[dishwasher_129]=True
    can_open[coffe_maker_130]=True
    can_open[microwave_135]=True
    can_open[window_191]=True
    can_open[nightstand_192]=True
    can_open[nightstand_195]=True
    can_open[bookshelf_196]=True
    can_open[filing_cabinet_200]=True
    can_open[curtain_204]=True
    can_open[curtain_205]=True
    can_open[curtain_206]=True
    can_open[dresser_274]=True
    can_open[bookshelf_275]=True
    can_open[curtain_289]=True
    can_open[curtain_290]=True
    can_open[curtain_291]=True
    can_open[window_310]=True
    can_open[diary_2008]=True
    can_open[envelope_2018]=True
    can_open[shampoo_2019]=True
    can_open[box_2038]=True
    can_open[pot_2040]=True
    can_open[after_shave_2042]=True
    can_open[stereo_2050]=True
    can_open[after_shave_2051]=True
    can_open[envelope_2055]=True
    can_open[tooth_paste_2059]=True
    can_open[novel_2060]=True
    can_open[after_shave_2063]=True
    has_switch[iron_2161]=True
    has_switch[washing_machine_2079]=True
    has_switch[remote_control_2124]=True
    has_switch[cd_player_2129]=True
    has_switch[dvd_player_2130]=True
    has_switch[stove_2135]=True
    has_switch[vacuum_cleaner_2139]=True
    has_switch[phone_2147]=True
    has_switch[faucet_20]=True
    has_switch[light_39]=True
    has_switch[phone_71]=True
    has_switch[light_73]=True
    has_switch[faucet_121]=True
    has_switch[fridge_126]=True
    has_switch[oven_127]=True
    has_switch[dishwasher_129]=True
    has_switch[coffe_maker_130]=True
    has_switch[toaster_132]=True
    has_switch[microwave_135]=True
    has_switch[computer_209]=True
    has_switch[light_212]=True
    has_switch[tablelamp_238]=True
    has_switch[tablelamp_239]=True
    has_switch[computer_276]=True
    has_switch[television_281]=True
    has_switch[light_283]=True
    has_switch[lighter_2004]=True
    has_switch[phone_2016]=True
    has_switch[phone_2017]=True
    has_switch[instrument_guitar_2028]=True
    has_switch[phone_2029]=True
    has_switch[laser_pointer_2034]=True
    has_switch[lighter_2039]=True
    has_switch[stereo_2050]=True
    has_switch[blow_dryer_2057]=True
    containers[basket_for_clothes_2078]=True
    containers[washing_machine_2079]=True
    containers[cd_player_2129]=True
    containers[stove_2135]=True
    containers[fryingpan_2154]=True
    containers[toilet_15]=True
    containers[bathroom_cabinet_17]=True
    containers[sink_19]=True
    containers[pot_78]=True
    containers[trashcan_99]=True
    containers[cupboard_117]=True
    containers[cupboard_118]=True
    containers[sink_120]=True
    containers[bookshelf_124]=True
    containers[fridge_126]=True
    containers[oven_127]=True
    containers[dishwasher_129]=True
    containers[coffe_maker_130]=True
    containers[toaster_132]=True
    containers[microwave_135]=True
    containers[nightstand_192]=True
    containers[nightstand_195]=True
    containers[bookshelf_196]=True
    containers[filing_cabinet_200]=True
    containers[dresser_274]=True
    containers[bookshelf_275]=True
    containers[box_2038]=True
    has_plug[iron_2161]=True
    has_plug[washing_machine_2079]=True
    has_plug[cd_player_2129]=True
    has_plug[dvd_player_2130]=True
    has_plug[vacuum_cleaner_2139]=True
    has_plug[phone_2147]=True
    has_plug[light_39]=True
    has_plug[phone_71]=True
    has_plug[light_73]=True
    has_plug[fridge_126]=True
    has_plug[oven_127]=True
    has_plug[coffe_maker_130]=True
    has_plug[toaster_132]=True
    has_plug[microwave_135]=True
    has_plug[keyboard_211]=True
    has_plug[light_212]=True
    has_plug[mouse_213]=True
    has_plug[keyboard_278]=True
    has_plug[mouse_280]=True
    has_plug[television_281]=True
    has_plug[light_283]=True
    has_plug[phone_2016]=True
    has_plug[phone_2017]=True
    has_plug[phone_2029]=True
    has_plug[stereo_2050]=True
    has_plug[blow_dryer_2057]=True
    readable[book_2136]=True
    readable[book_2137]=True
    readable[diary_2008]=True
    readable[check_2026]=True
    readable[homework_2047]=True
    readable[check_2058]=True
    readable[novel_2060]=True
    readable[check_2071]=True
    readable[check_2075]=True
    lookable[drawing_33]=True
    lookable[drawing_110]=True
    lookable[drawing_111]=True
    lookable[drawing_201]=True
    lookable[drawing_202]=True
    lookable[computer_209]=True
    lookable[computer_276]=True
    lookable[television_281]=True
    lookable[drawing_288]=True
    is_clothes[clothes_pants_2157]=True
    is_clothes[clothes_shirt_2158]=True
    is_clothes[clothes_socks_2159]=True
    is_clothes[clothes_skirt_2160]=True
    is_clothes[clothes_dress_2116]=True
    is_clothes[clothes_hat_2117]=True
    is_clothes[clothes_gloves_2118]=True
    is_clothes[clothes_jacket_2119]=True
    is_clothes[clothes_scarf_2120]=True
    is_clothes[clothes_underwear_2121]=True
    is_clothes[headset_2131]=True
    is_clothes[headset_2146]=True
    is_clothes[spectacles_2153]=True
    is_clothes[shoes_2033]=True
    is_clothes[clothes_pants_2036]=True
    is_food[food_steak_2080]=True
    is_food[food_apple_2081]=True
    is_food[food_bacon_2082]=True
    is_food[food_banana_2083]=True
    is_food[food_bread_2084]=True
    is_food[food_cake_2085]=True
    is_food[food_carrot_2086]=True
    is_food[food_cereal_2087]=True
    is_food[food_cheese_2088]=True
    is_food[food_chicken_2089]=True
    is_food[food_dessert_2090]=True
    is_food[food_donut_2091]=True
    is_food[food_egg_2092]=True
    is_food[food_fish_2093]=True
    is_food[food_food_2094]=True
    is_food[food_fruit_2095]=True
    is_food[food_hamburger_2096]=True
    is_food[food_ice_cream_2097]=True
    is_food[food_jam_2098]=True
    is_food[food_kiwi_2099]=True
    is_food[food_lemon_2100]=True
    is_food[food_noodles_2101]=True
    is_food[food_oatmeal_2102]=True
    is_food[food_orange_2103]=True
    is_food[food_onion_2104]=True
    is_food[food_peanut_butter_2105]=True
    is_food[food_pizza_2106]=True
    is_food[food_potato_2107]=True
    is_food[food_rice_2108]=True
    is_food[food_salt_2109]=True
    is_food[food_snack_2110]=True
    is_food[food_sugar_2111]=True
    is_food[food_turkey_2112]=True
    is_food[food_vegetable_2113]=True
    is_food[food_food_1000]=True
    is_food[food_food_2001]=True
    is_food[food_butter_2007]=True
    is_food[food_onion_2009]=True
    is_food[food_carrot_2015]=True
    is_food[food_food_2021]=True
    is_food[food_orange_2027]=True
    is_food[food_salt_2041]=True
    is_food[food_food_2046]=True
    is_food[food_onion_2048]=True
    is_food[food_kiwi_2054]=True
    is_food[food_orange_2061]=True
    is_food[food_food_2064]=True
    is_food[food_cheese_2072]=True
    is_food[food_food_2073]=True
    is_food[food_food_2074]=True
    is_food[food_peanut_butter_2077]=True
    cover_object[towel_2128]=True
    cover_object[curtain_22]=True
    cover_object[curtain_204]=True
    cover_object[curtain_205]=True
    cover_object[curtain_206]=True
    cover_object[curtain_289]=True
    cover_object[curtain_290]=True
    cover_object[curtain_291]=True
    cover_object[table_cloth_2005]=True
    cover_object[envelope_2018]=True
    cover_object[rag_2025]=True
    cover_object[box_2038]=True
    cover_object[rag_2052]=True
    cover_object[envelope_2055]=True
    cover_object[toilet_paper_2076]=True
    has_paper[book_2136]=True
    has_paper[book_2137]=True
    has_paper[drawing_33]=True
    has_paper[drawing_110]=True
    has_paper[drawing_111]=True
    has_paper[drawing_201]=True
    has_paper[drawing_202]=True
    has_paper[drawing_288]=True
    has_paper[diary_2008]=True
    has_paper[envelope_2018]=True
    has_paper[check_2026]=True
    has_paper[homework_2047]=True
    has_paper[coffee_filter_2053]=True
    has_paper[envelope_2055]=True
    has_paper[check_2058]=True
    has_paper[novel_2060]=True
    has_paper[coffee_filter_2065]=True
    has_paper[check_2071]=True
    has_paper[check_2075]=True
    has_paper[toilet_paper_2076]=True
    movable[clothes_pants_2157]=True
    movable[clothes_shirt_2158]=True
    movable[clothes_socks_2159]=True
    movable[clothes_skirt_2160]=True
    movable[iron_2161]=True
    movable[basket_for_clothes_2078]=True
    movable[food_steak_2080]=True
    movable[food_apple_2081]=True
    movable[food_bacon_2082]=True
    movable[food_banana_2083]=True
    movable[food_bread_2084]=True
    movable[food_cake_2085]=True
    movable[food_carrot_2086]=True
    movable[food_cereal_2087]=True
    movable[food_cheese_2088]=True
    movable[food_chicken_2089]=True
    movable[food_dessert_2090]=True
    movable[food_donut_2091]=True
    movable[food_egg_2092]=True
    movable[food_fish_2093]=True
    movable[food_food_2094]=True
    movable[food_fruit_2095]=True
    movable[food_hamburger_2096]=True
    movable[food_ice_cream_2097]=True
    movable[food_jam_2098]=True
    movable[food_kiwi_2099]=True
    movable[food_lemon_2100]=True
    movable[food_noodles_2101]=True
    movable[food_oatmeal_2102]=True
    movable[food_orange_2103]=True
    movable[food_onion_2104]=True
    movable[food_peanut_butter_2105]=True
    movable[food_pizza_2106]=True
    movable[food_potato_2107]=True
    movable[food_rice_2108]=True
    movable[food_salt_2109]=True
    movable[food_snack_2110]=True
    movable[food_sugar_2111]=True
    movable[food_turkey_2112]=True
    movable[food_vegetable_2113]=True
    movable[dry_pasta_2114]=True
    movable[milk_2115]=True
    movable[clothes_dress_2116]=True
    movable[clothes_hat_2117]=True
    movable[clothes_gloves_2118]=True
    movable[clothes_jacket_2119]=True
    movable[clothes_scarf_2120]=True
    movable[clothes_underwear_2121]=True
    movable[knife_2122]=True
    movable[cutting_board_2123]=True
    movable[remote_control_2124]=True
    movable[soap_2125]=True
    movable[soap_2126]=True
    movable[towel_2128]=True
    movable[cd_player_2129]=True
    movable[dvd_player_2130]=True
    movable[headset_2131]=True
    movable[cup_2132]=True
    movable[cup_2133]=True
    movable[cup_2134]=True
    movable[book_2136]=True
    movable[book_2137]=True
    movable[pot_2138]=True
    movable[vacuum_cleaner_2139]=True
    movable[bowl_2140]=True
    movable[bowl_2141]=True
    movable[bowl_2142]=True
    movable[cleaning_solution_2143]=True
    movable[ironing_board_2144]=True
    movable[cd_2145]=True
    movable[headset_2146]=True
    movable[phone_2147]=True
    movable[sauce_2148]=True
    movable[oil_2149]=True
    movable[fork_2150]=True
    movable[fork_2151]=True
    movable[plate_2152]=True
    movable[spectacles_2153]=True
    movable[fryingpan_2154]=True
    movable[detergent_2155]=True
    movable[curtain_22]=True
    movable[mat_32]=True
    movable[drawing_33]=True
    movable[phone_71]=True
    movable[pot_78]=True
    movable[trashcan_99]=True
    movable[mat_102]=True
    movable[pillow_103]=True
    movable[pillow_104]=True
    movable[pillow_105]=True
    movable[pillow_106]=True
    movable[pillow_107]=True
    movable[pillow_108]=True
    movable[drawing_110]=True
    movable[drawing_111]=True
    movable[bench_113]=True
    movable[table_114]=True
    movable[bench_115]=True
    movable[tray_128]=True
    movable[coffe_maker_130]=True
    movable[toaster_132]=True
    movable[desk_193]=True
    movable[chair_194]=True
    movable[couch_198]=True
    movable[table_199]=True
    movable[drawing_201]=True
    movable[drawing_202]=True
    movable[mat_203]=True
    movable[curtain_204]=True
    movable[curtain_205]=True
    movable[curtain_206]=True
    movable[pillow_207]=True
    movable[pillow_208]=True
    movable[keyboard_211]=True
    movable[mouse_213]=True
    movable[mousepad_214]=True
    movable[couch_269]=True
    movable[table_270]=True
    movable[chair_271]=True
    movable[desk_272]=True
    movable[keyboard_278]=True
    movable[mousepad_279]=True
    movable[mouse_280]=True
    movable[mat_284]=True
    movable[pillow_286]=True
    movable[pillow_287]=True
    movable[drawing_288]=True
    movable[curtain_289]=True
    movable[curtain_290]=True
    movable[curtain_291]=True
    movable[hanger_292]=True
    movable[hanger_293]=True
    movable[hanger_294]=True
    movable[food_food_1000]=True
    movable[wooden_spoon_2000]=True
    movable[food_food_2001]=True
    movable[brush_2002]=True
    movable[chair_2003]=True
    movable[lighter_2004]=True
    movable[table_cloth_2005]=True
    movable[piano_bench_2006]=True
    movable[food_butter_2007]=True
    movable[diary_2008]=True
    movable[food_onion_2009]=True
    movable[soap_2010]=True
    movable[detergent_2011]=True
    movable[measuring_cup_2012]=True
    movable[oil_2013]=True
    movable[pencil_2014]=True
    movable[food_carrot_2015]=True
    movable[phone_2016]=True
    movable[phone_2017]=True
    movable[envelope_2018]=True
    movable[shampoo_2019]=True
    movable[pencil_2020]=True
    movable[food_food_2021]=True
    movable[stamp_2022]=True
    movable[tea_bag_2023]=True
    movable[ice_2024]=True
    movable[rag_2025]=True
    movable[check_2026]=True
    movable[food_orange_2027]=True
    movable[instrument_guitar_2028]=True
    movable[phone_2029]=True
    movable[cd_2030]=True
    movable[scrabble_2031]=True
    movable[shoes_2033]=True
    movable[laser_pointer_2034]=True
    movable[knife_2035]=True
    movable[clothes_pants_2036]=True
    movable[knife_2037]=True
    movable[box_2038]=True
    movable[lighter_2039]=True
    movable[pot_2040]=True
    movable[food_salt_2041]=True
    movable[after_shave_2042]=True
    movable[stamp_2043]=True
    movable[shoe_rack_2044]=True
    movable[glue_2045]=True
    movable[food_food_2046]=True
    movable[homework_2047]=True
    movable[food_onion_2048]=True
    movable[cup_2049]=True
    movable[stereo_2050]=True
    movable[after_shave_2051]=True
    movable[rag_2052]=True
    movable[coffee_filter_2053]=True
    movable[food_kiwi_2054]=True
    movable[envelope_2055]=True
    movable[toy_2056]=True
    movable[blow_dryer_2057]=True
    movable[check_2058]=True
    movable[tooth_paste_2059]=True
    movable[novel_2060]=True
    movable[food_orange_2061]=True
    movable[piano_bench_2062]=True
    movable[after_shave_2063]=True
    movable[food_food_2064]=True
    movable[coffee_filter_2065]=True
    movable[tea_2066]=True
    movable[piano_bench_2067]=True
    movable[tray_2068]=True
    movable[cat_2069]=True
    movable[chessboard_2070]=True
    movable[check_2071]=True
    movable[food_cheese_2072]=True
    movable[food_food_2073]=True
    movable[food_food_2074]=True
    movable[check_2075]=True
    movable[toilet_paper_2076]=True
    movable[food_peanut_butter_2077]=True
    cream[food_cheese_2088]=True
    cream[food_ice_cream_2097]=True
    cream[food_jam_2098]=True
    cream[food_peanut_butter_2105]=True
    cream[soap_2125]=True
    cream[soap_2126]=True
    cream[sauce_2148]=True
    cream[food_butter_2007]=True
    cream[soap_2010]=True
    cream[after_shave_2042]=True
    cream[glue_2045]=True
    cream[after_shave_2051]=True
    cream[tooth_paste_2059]=True
    cream[after_shave_2063]=True
    cream[food_cheese_2072]=True
    cream[food_peanut_butter_2077]=True
    #properties_end

    #relations
    on[iron_2161,bowl_2142]=True
    on[clothes_dress_2116,bed_197]=True
    on[clothes_hat_2117,table_114]=True
    on[clothes_gloves_2118,table_114]=True
    on[clothes_jacket_2119,couch_198]=True
    on[knife_2122,table_114]=True
    on[cutting_board_2123,kitchen_counter_119]=True
    on[remote_control_2124,tvstand_273]=True
    on[soap_2125,sink_19]=True
    on[soap_2126,sink_120]=True
    on[cd_player_2129,tvstand_273]=True
    on[dvd_player_2130,tvstand_273]=True
    on[headset_2131,tvstand_273]=True
    on[cup_2132,table_114]=True
    on[cup_2133,table_114]=True
    on[cup_2134,table_114]=True
    on[stove_2135,kitchen_counter_119]=True
    on[book_2136,bookshelf_124]=True
    on[book_2137,bookshelf_124]=True
    on[pot_2138,kitchen_counter_119]=True
    on[bowl_2140,kitchen_counter_119]=True
    on[bowl_2141,kitchen_counter_119]=True
    on[bowl_2142,kitchen_counter_119]=True
    on[cleaning_solution_2143,sink_19]=True
    on[cd_2145,tvstand_273]=True
    on[headset_2146,desk_272]=True
    on[phone_2147,desk_272]=True
    on[oil_2149,kitchen_counter_123]=True
    on[fork_2150,kitchen_counter_119]=True
    on[fork_2151,kitchen_counter_119]=True
    on[plate_2152,kitchen_counter_119]=True
    on[spectacles_2153,kitchen_counter_122]=True
    on[fryingpan_2154,kitchen_counter_122]=True
    on[detergent_2155,sink_19]=True
    on[ceiling_6,wall_3]=True
    on[ceiling_7,wall_2]=True
    on[ceiling_8,wall_5]=True
    on[ceiling_9,wall_4]=True
    on[faucet_20,bathroom_counter_18]=True
    on[shower_21,floor_13]=True
    on[door_38,floor_12]=True
    on[ceiling_52,wall_70]=True
    on[ceiling_54,wall_67]=True
    on[ceiling_58,wall_69]=True
    on[ceiling_60,wall_68]=True
    on[door_61,floor_169]=True
    on[door_62,floor_261]=True
    on[knifeblock_76,wall_64]=True
    on[pot_78,oven_127]=True
    on[trashcan_99,floor_51]=True
    on[mat_102,floor_47]=True
    on[pillow_103,bench_113]=True
    on[pillow_104,bench_113]=True
    on[pillow_105,bench_115]=True
    on[pillow_106,bench_115]=True
    on[pillow_107,tvstand_116]=True
    on[pillow_108,tvstand_116]=True
    on[drawing_110,bookshelf_124]=True
    on[table_114,floor_47]=True
    on[table_114,mat_102]=True
    on[tvstand_116,floor_48]=True
    on[cupboard_117,wall_67]=True
    on[cupboard_118,wall_68]=True
    on[faucet_121,kitchen_counter_119]=True
    on[kitchen_counter_123,floor_45]=True
    on[bookshelf_124,floor_42]=True
    on[bookshelf_124,floor_43]=True
    on[fridge_126,floor_44]=True
    on[coffe_maker_130,kitchen_counter_122]=True
    on[toaster_132,kitchen_counter_122]=True
    on[microwave_135,kitchen_counter_122]=True
    on[ceiling_181,wall_175]=True
    on[ceiling_183,wall_176]=True
    on[ceiling_187,wall_178]=True
    on[ceiling_189,wall_177]=True
    on[nightstand_192,floor_166]=True
    on[desk_193,floor_163]=True
    on[desk_193,floor_164]=True
    on[nightstand_195,floor_165]=True
    on[bookshelf_196,floor_170]=True
    on[filing_cabinet_200,floor_170]=True
    on[pillow_207,bed_197]=True
    on[pillow_208,bed_197]=True
    on[cpuscreen_210,desk_193]=True
    on[keyboard_211,desk_193]=True
    on[mouse_213,desk_193]=True
    on[mouse_213,mousepad_214]=True
    on[mousepad_214,desk_193]=True
    on[tablelamp_238,nightstand_192]=True
    on[tablelamp_239,nightstand_195]=True
    on[ceiling_250,wall_247]=True
    on[ceiling_252,wall_246]=True
    on[ceiling_256,wall_248]=True
    on[ceiling_258,wall_249]=True
    on[desk_272,floor_263]=True
    on[tvstand_273,floor_259]=True
    on[tvstand_273,floor_260]=True
    on[bookshelf_275,floor_262]=True
    on[cpuscreen_277,desk_272]=True
    on[keyboard_278,desk_272]=True
    on[mousepad_279,desk_272]=True
    on[mouse_280,desk_272]=True
    on[mouse_280,mousepad_279]=True
    on[television_281,tvstand_273]=True
    on[orchid_285,table_270]=True
    on[curtain_291,couch_269]=True
    on[wooden_spoon_2000,table_199]=True
    on[brush_2002,couch_269]=True
    on[chair_2003,couch_198]=True
    on[lighter_2004,mat_102]=True
    on[table_cloth_2005,table_114]=True
    on[piano_bench_2006,floor_44]=True
    on[food_butter_2007,table_cloth_2005]=True
    on[pencil_2014,table_270]=True
    on[phone_2016,couch_198]=True
    on[phone_2017,couch_269]=True
    on[shampoo_2019,table_270]=True
    on[pencil_2020,bookshelf_275]=True
    on[food_food_2021,table_114]=True
    on[stamp_2022,desk_272]=True
    on[tea_bag_2023,table_199]=True
    on[check_2026,desk_193]=True
    on[food_orange_2027,kitchen_counter_123]=True
    on[instrument_guitar_2028,couch_198]=True
    on[phone_2029,bathroom_counter_18]=True
    on[shoes_2033,couch_269]=True
    on[laser_pointer_2034,desk_193]=True
    on[knife_2035,kitchen_counter_123]=True
    on[clothes_pants_2036,hanger_292]=True
    on[box_2038,table_114]=True
    on[lighter_2039,mat_102]=True
    on[food_salt_2041,kitchen_counter_119]=True
    on[stamp_2043,desk_272]=True
    on[shoe_rack_2044,mat_203]=True
    on[cup_2049,table_114]=True
    on[rag_2052,couch_198]=True
    on[food_kiwi_2054,kitchen_counter_123]=True
    on[envelope_2055,bookshelf_124]=True
    on[toy_2056,mat_32]=True
    on[check_2058,table_114]=True
    on[novel_2060,bookshelf_196]=True
    on[piano_bench_2062,floor_44]=True
    on[food_food_2064,oven_127]=True
    on[piano_bench_2067,mat_32]=True
    on[tray_2068,kitchen_counter_123]=True
    on[chessboard_2070,shoe_rack_2044]=True
    on[check_2071,shoe_rack_2044]=True
    inside[clothes_pants_2157,basket_for_clothes_2078]=True
    inside[clothes_pants_2157,dining_room_41]=True
    inside[clothes_shirt_2158,basket_for_clothes_2078]=True
    inside[clothes_shirt_2158,dining_room_41]=True
    inside[clothes_socks_2159,basket_for_clothes_2078]=True
    inside[clothes_socks_2159,dining_room_41]=True
    inside[clothes_skirt_2160,basket_for_clothes_2078]=True
    inside[clothes_skirt_2160,dining_room_41]=True
    inside[iron_2161,dining_room_41]=True
    inside[basket_for_clothes_2078,dining_room_41]=True
    inside[washing_machine_2079,dining_room_41]=True
    inside[food_steak_2080,dining_room_41]=True
    inside[food_steak_2080,fridge_126]=True
    inside[food_apple_2081,dining_room_41]=True
    inside[food_apple_2081,fridge_126]=True
    inside[food_bacon_2082,dining_room_41]=True
    inside[food_bacon_2082,fridge_126]=True
    inside[food_banana_2083,dining_room_41]=True
    inside[food_banana_2083,fridge_126]=True
    inside[food_bread_2084,dining_room_41]=True
    inside[food_bread_2084,table_114]=True
    inside[food_cake_2085,dining_room_41]=True
    inside[food_cake_2085,fridge_126]=True
    inside[food_carrot_2086,dining_room_41]=True
    inside[food_carrot_2086,fridge_126]=True
    inside[food_cereal_2087,dining_room_41]=True
    inside[food_cereal_2087,fridge_126]=True
    inside[food_cheese_2088,dining_room_41]=True
    inside[food_cheese_2088,fridge_126]=True
    inside[food_chicken_2089,dining_room_41]=True
    inside[food_chicken_2089,fridge_126]=True
    inside[food_dessert_2090,dining_room_41]=True
    inside[food_dessert_2090,fridge_126]=True
    inside[food_donut_2091,dining_room_41]=True
    inside[food_donut_2091,fridge_126]=True
    inside[food_egg_2092,dining_room_41]=True
    inside[food_egg_2092,fridge_126]=True
    inside[food_fish_2093,dining_room_41]=True
    inside[food_fish_2093,fridge_126]=True
    inside[food_food_2094,dining_room_41]=True
    inside[food_food_2094,fridge_126]=True
    inside[food_fruit_2095,dining_room_41]=True
    inside[food_fruit_2095,fridge_126]=True
    inside[food_hamburger_2096,dining_room_41]=True
    inside[food_hamburger_2096,fridge_126]=True
    inside[food_ice_cream_2097,dining_room_41]=True
    inside[food_ice_cream_2097,fridge_126]=True
    inside[food_jam_2098,dining_room_41]=True
    inside[food_jam_2098,fridge_126]=True
    inside[food_kiwi_2099,dining_room_41]=True
    inside[food_kiwi_2099,fridge_126]=True
    inside[food_lemon_2100,dining_room_41]=True
    inside[food_lemon_2100,fridge_126]=True
    inside[food_noodles_2101,dining_room_41]=True
    inside[food_noodles_2101,fridge_126]=True
    inside[food_oatmeal_2102,dining_room_41]=True
    inside[food_oatmeal_2102,fridge_126]=True
    inside[food_orange_2103,dining_room_41]=True
    inside[food_orange_2103,fridge_126]=True
    inside[food_onion_2104,dining_room_41]=True
    inside[food_onion_2104,fridge_126]=True
    inside[food_peanut_butter_2105,dining_room_41]=True
    inside[food_peanut_butter_2105,fridge_126]=True
    inside[food_pizza_2106,dining_room_41]=True
    inside[food_pizza_2106,fridge_126]=True
    inside[food_potato_2107,dining_room_41]=True
    inside[food_potato_2107,fridge_126]=True
    inside[food_rice_2108,dining_room_41]=True
    inside[food_rice_2108,fridge_126]=True
    inside[food_salt_2109,dining_room_41]=True
    inside[food_salt_2109,fridge_126]=True
    inside[food_snack_2110,dining_room_41]=True
    inside[food_snack_2110,fridge_126]=True
    inside[food_sugar_2111,dining_room_41]=True
    inside[food_sugar_2111,fridge_126]=True
    inside[food_turkey_2112,dining_room_41]=True
    inside[food_turkey_2112,fridge_126]=True
    inside[food_vegetable_2113,dining_room_41]=True
    inside[food_vegetable_2113,fridge_126]=True
    inside[dry_pasta_2114,dining_room_41]=True
    inside[dry_pasta_2114,table_114]=True
    inside[milk_2115,dining_room_41]=True
    inside[milk_2115,table_114]=True
    inside[clothes_dress_2116,bedroom_162]=True
    inside[clothes_hat_2117,dining_room_41]=True
    inside[clothes_gloves_2118,dining_room_41]=True
    inside[clothes_jacket_2119,bedroom_162]=True
    inside[clothes_scarf_2120,bedroom_162]=True
    inside[clothes_scarf_2120,bed_197]=True
    inside[clothes_underwear_2121,bedroom_162]=True
    inside[clothes_underwear_2121,bed_197]=True
    inside[knife_2122,dining_room_41]=True
    inside[cutting_board_2123,dining_room_41]=True
    inside[remote_control_2124,home_office_241]=True
    inside[soap_2125,bathroom_1]=True
    inside[soap_2126,dining_room_41]=True
    inside[towel_2128,bathroom_1]=True
    inside[towel_2128,drawing_33]=True
    inside[cd_player_2129,home_office_241]=True
    inside[dvd_player_2130,home_office_241]=True
    inside[headset_2131,home_office_241]=True
    inside[cup_2132,dining_room_41]=True
    inside[cup_2133,dining_room_41]=True
    inside[cup_2134,dining_room_41]=True
    inside[stove_2135,dining_room_41]=True
    inside[book_2136,dining_room_41]=True
    inside[book_2137,dining_room_41]=True
    inside[pot_2138,dining_room_41]=True
    inside[vacuum_cleaner_2139,dining_room_41]=True
    inside[bowl_2140,dining_room_41]=True
    inside[bowl_2141,dining_room_41]=True
    inside[bowl_2142,dining_room_41]=True
    inside[cleaning_solution_2143,bathroom_1]=True
    inside[ironing_board_2144,dining_room_41]=True
    inside[cd_2145,home_office_241]=True
    inside[headset_2146,home_office_241]=True
    inside[phone_2147,home_office_241]=True
    inside[sauce_2148,dining_room_41]=True
    inside[sauce_2148,fridge_126]=True
    inside[oil_2149,dining_room_41]=True
    inside[fork_2150,dining_room_41]=True
    inside[fork_2151,dining_room_41]=True
    inside[plate_2152,dining_room_41]=True
    inside[spectacles_2153,dining_room_41]=True
    inside[fryingpan_2154,dining_room_41]=True
    inside[detergent_2155,bathroom_1]=True
    inside[window_2156,bathroom_1]=True
    inside[wall_2,bathroom_1]=True
    inside[wall_3,bathroom_1]=True
    inside[wall_4,bathroom_1]=True
    inside[wall_5,bathroom_1]=True
    inside[ceiling_6,bathroom_1]=True
    inside[ceiling_7,bathroom_1]=True
    inside[ceiling_8,bathroom_1]=True
    inside[ceiling_9,bathroom_1]=True
    inside[floor_10,bathroom_1]=True
    inside[floor_11,bathroom_1]=True
    inside[floor_12,bathroom_1]=True
    inside[floor_13,bathroom_1]=True
    inside[floor_14,bathroom_1]=True
    inside[toilet_15,bathroom_1]=True
    inside[shower_16,bathroom_1]=True
    inside[bathroom_cabinet_17,bathroom_1]=True
    inside[bathroom_counter_18,bathroom_1]=True
    inside[sink_19,bathroom_1]=True
    inside[sink_19,bathroom_counter_18]=True
    inside[faucet_20,bathroom_1]=True
    inside[shower_21,bathroom_1]=True
    inside[curtain_22,bathroom_1]=True
    inside[curtain_22,shower_21]=True
    inside[mat_32,bathroom_1]=True
    inside[drawing_33,bathroom_1]=True
    inside[walllamp_34,bathroom_1]=True
    inside[ceilinglamp_35,bathroom_1]=True
    inside[walllamp_36,bathroom_1]=True
    inside[doorjamb_37,bathroom_1]=True
    inside[door_38,bathroom_1]=True
    inside[light_39,bathroom_1]=True
    inside[floor_42,dining_room_41]=True
    inside[floor_43,dining_room_41]=True
    inside[floor_44,dining_room_41]=True
    inside[floor_45,dining_room_41]=True
    inside[floor_46,dining_room_41]=True
    inside[floor_47,dining_room_41]=True
    inside[floor_48,dining_room_41]=True
    inside[floor_49,dining_room_41]=True
    inside[floor_50,dining_room_41]=True
    inside[floor_51,dining_room_41]=True
    inside[ceiling_52,dining_room_41]=True
    inside[ceiling_53,dining_room_41]=True
    inside[ceiling_54,dining_room_41]=True
    inside[ceiling_55,dining_room_41]=True
    inside[ceiling_56,dining_room_41]=True
    inside[ceiling_57,dining_room_41]=True
    inside[ceiling_58,dining_room_41]=True
    inside[ceiling_59,dining_room_41]=True
    inside[ceiling_60,dining_room_41]=True
    inside[door_61,dining_room_41]=True
    inside[door_62,dining_room_41]=True
    inside[wall_63,dining_room_41]=True
    inside[wall_64,dining_room_41]=True
    inside[wall_65,dining_room_41]=True
    inside[wall_66,dining_room_41]=True
    inside[wall_67,dining_room_41]=True
    inside[wall_68,dining_room_41]=True
    inside[wall_69,dining_room_41]=True
    inside[wall_70,dining_room_41]=True
    inside[phone_71,dining_room_41]=True
    inside[powersocket_72,dining_room_41]=True
    inside[light_73,dining_room_41]=True
    inside[knifeblock_76,dining_room_41]=True
    inside[pot_78,dining_room_41]=True
    inside[trashcan_99,dining_room_41]=True
    inside[mat_102,dining_room_41]=True
    inside[pillow_103,dining_room_41]=True
    inside[pillow_104,dining_room_41]=True
    inside[pillow_105,dining_room_41]=True
    inside[pillow_106,dining_room_41]=True
    inside[pillow_107,dining_room_41]=True
    inside[pillow_108,dining_room_41]=True
    inside[drawing_110,dining_room_41]=True
    inside[drawing_111,dining_room_41]=True
    inside[bench_113,dining_room_41]=True
    inside[table_114,dining_room_41]=True
    inside[bench_115,dining_room_41]=True
    inside[tvstand_116,dining_room_41]=True
    inside[cupboard_117,dining_room_41]=True
    inside[cupboard_118,dining_room_41]=True
    inside[kitchen_counter_119,dining_room_41]=True
    inside[sink_120,dining_room_41]=True
    inside[sink_120,kitchen_counter_119]=True
    inside[faucet_121,dining_room_41]=True
    inside[kitchen_counter_122,dining_room_41]=True
    inside[kitchen_counter_123,dining_room_41]=True
    inside[bookshelf_124,dining_room_41]=True
    inside[stovefan_125,dining_room_41]=True
    inside[fridge_126,dining_room_41]=True
    inside[oven_127,dining_room_41]=True
    inside[tray_128,dining_room_41]=True
    inside[tray_128,oven_127]=True
    inside[dishwasher_129,dining_room_41]=True
    inside[coffe_maker_130,dining_room_41]=True
    inside[toaster_132,dining_room_41]=True
    inside[microwave_135,dining_room_41]=True
    inside[ceilinglamp_137,dining_room_41]=True
    inside[ceilinglamp_138,dining_room_41]=True
    inside[walllamp_139,dining_room_41]=True
    inside[walllamp_140,dining_room_41]=True
    inside[walllamp_141,dining_room_41]=True
    inside[floor_163,bedroom_162]=True
    inside[floor_164,bedroom_162]=True
    inside[floor_165,bedroom_162]=True
    inside[floor_166,bedroom_162]=True
    inside[floor_167,bedroom_162]=True
    inside[floor_168,bedroom_162]=True
    inside[floor_169,bedroom_162]=True
    inside[floor_170,bedroom_162]=True
    inside[floor_171,bedroom_162]=True
    inside[floor_172,bedroom_162]=True
    inside[wall_173,bedroom_162]=True
    inside[wall_174,bedroom_162]=True
    inside[wall_175,bedroom_162]=True
    inside[wall_176,bedroom_162]=True
    inside[wall_177,bedroom_162]=True
    inside[wall_178,bedroom_162]=True
    inside[wall_179,bedroom_162]=True
    inside[wall_180,bedroom_162]=True
    inside[ceiling_181,bedroom_162]=True
    inside[ceiling_182,bedroom_162]=True
    inside[ceiling_183,bedroom_162]=True
    inside[ceiling_184,bedroom_162]=True
    inside[ceiling_185,bedroom_162]=True
    inside[ceiling_186,bedroom_162]=True
    inside[ceiling_187,bedroom_162]=True
    inside[ceiling_188,bedroom_162]=True
    inside[ceiling_189,bedroom_162]=True
    inside[doorjamb_190,bedroom_162]=True
    inside[window_191,bedroom_162]=True
    inside[nightstand_192,bedroom_162]=True
    inside[desk_193,bedroom_162]=True
    inside[chair_194,bedroom_162]=True
    inside[nightstand_195,bedroom_162]=True
    inside[bookshelf_196,bedroom_162]=True
    inside[bed_197,bedroom_162]=True
    inside[couch_198,bedroom_162]=True
    inside[table_199,bedroom_162]=True
    inside[filing_cabinet_200,bedroom_162]=True
    inside[drawing_201,bedroom_162]=True
    inside[drawing_202,bedroom_162]=True
    inside[mat_203,bedroom_162]=True
    inside[curtain_204,bedroom_162]=True
    inside[curtain_204,curtain_205]=True
    inside[curtain_205,bedroom_162]=True
    inside[curtain_205,curtain_204]=True
    inside[curtain_206,bedroom_162]=True
    inside[pillow_207,bedroom_162]=True
    inside[pillow_208,bedroom_162]=True
    inside[computer_209,bedroom_162]=True
    inside[cpuscreen_210,bedroom_162]=True
    inside[keyboard_211,bedroom_162]=True
    inside[light_212,bedroom_162]=True
    inside[mouse_213,bedroom_162]=True
    inside[mousepad_214,bedroom_162]=True
    inside[photoframe_219,bedroom_162]=True
    inside[photoframe_219,bookshelf_196]=True
    inside[ceilinglamp_237,bedroom_162]=True
    inside[tablelamp_238,bedroom_162]=True
    inside[tablelamp_239,bedroom_162]=True
    inside[wall_242,home_office_241]=True
    inside[wall_243,home_office_241]=True
    inside[wall_244,home_office_241]=True
    inside[wall_245,home_office_241]=True
    inside[wall_246,home_office_241]=True
    inside[wall_247,home_office_241]=True
    inside[wall_248,home_office_241]=True
    inside[wall_249,home_office_241]=True
    inside[ceiling_250,home_office_241]=True
    inside[ceiling_251,home_office_241]=True
    inside[ceiling_252,home_office_241]=True
    inside[ceiling_253,home_office_241]=True
    inside[ceiling_254,home_office_241]=True
    inside[ceiling_255,home_office_241]=True
    inside[ceiling_256,home_office_241]=True
    inside[ceiling_257,home_office_241]=True
    inside[ceiling_258,home_office_241]=True
    inside[floor_259,home_office_241]=True
    inside[floor_260,home_office_241]=True
    inside[floor_261,home_office_241]=True
    inside[floor_262,home_office_241]=True
    inside[floor_263,home_office_241]=True
    inside[floor_264,home_office_241]=True
    inside[floor_265,home_office_241]=True
    inside[floor_266,home_office_241]=True
    inside[floor_267,home_office_241]=True
    inside[floor_268,home_office_241]=True
    inside[couch_269,home_office_241]=True
    inside[table_270,home_office_241]=True
    inside[table_270,couch_269]=True
    inside[chair_271,home_office_241]=True
    inside[desk_272,home_office_241]=True
    inside[tvstand_273,home_office_241]=True
    inside[dresser_274,home_office_241]=True
    inside[bookshelf_275,home_office_241]=True
    inside[computer_276,home_office_241]=True
    inside[cpuscreen_277,home_office_241]=True
    inside[keyboard_278,home_office_241]=True
    inside[mousepad_279,home_office_241]=True
    inside[mouse_280,home_office_241]=True
    inside[television_281,home_office_241]=True
    inside[powersocket_282,home_office_241]=True
    inside[light_283,home_office_241]=True
    inside[mat_284,home_office_241]=True
    inside[orchid_285,home_office_241]=True
    inside[orchid_285,couch_269]=True
    inside[pillow_286,home_office_241]=True
    inside[pillow_286,couch_269]=True
    inside[pillow_287,home_office_241]=True
    inside[pillow_287,couch_269]=True
    inside[drawing_288,home_office_241]=True
    inside[curtain_289,home_office_241]=True
    inside[curtain_289,curtain_290]=True
    inside[curtain_290,home_office_241]=True
    inside[curtain_290,curtain_289]=True
    inside[curtain_291,home_office_241]=True
    inside[hanger_292,home_office_241]=True
    inside[hanger_292,dresser_274]=True
    inside[hanger_293,home_office_241]=True
    inside[hanger_293,dresser_274]=True
    inside[hanger_294,home_office_241]=True
    inside[hanger_294,dresser_274]=True
    inside[ceilinglamp_303,home_office_241]=True
    inside[walllamp_304,home_office_241]=True
    inside[walllamp_305,home_office_241]=True
    inside[walllamp_306,home_office_241]=True
    inside[walllamp_307,home_office_241]=True
    inside[doorjamb_309,home_office_241]=True
    inside[window_310,home_office_241]=True
    inside[food_food_1000,dining_room_41]=True
    inside[wooden_spoon_2000,bedroom_162]=True
    inside[food_food_2001,dining_room_41]=True
    inside[food_food_2001,fridge_126]=True
    inside[brush_2002,home_office_241]=True
    inside[chair_2003,bedroom_162]=True
    inside[lighter_2004,dining_room_41]=True
    inside[table_cloth_2005,dining_room_41]=True
    inside[piano_bench_2006,dining_room_41]=True
    inside[food_butter_2007,dining_room_41]=True
    inside[diary_2008,bedroom_162]=True
    inside[diary_2008,filing_cabinet_200]=True
    inside[food_onion_2009,dining_room_41]=True
    inside[food_onion_2009,trashcan_99]=True
    inside[soap_2010,dining_room_41]=True
    inside[soap_2010,sink_120]=True
    inside[detergent_2011,dining_room_41]=True
    inside[detergent_2011,dishwasher_129]=True
    inside[measuring_cup_2012,dining_room_41]=True
    inside[measuring_cup_2012,dishwasher_129]=True
    inside[oil_2013,dining_room_41]=True
    inside[oil_2013,oven_127]=True
    inside[pencil_2014,home_office_241]=True
    inside[food_carrot_2015,dining_room_41]=True
    inside[food_carrot_2015,oven_127]=True
    inside[phone_2016,bedroom_162]=True
    inside[phone_2017,home_office_241]=True
    inside[envelope_2018,bedroom_162]=True
    inside[envelope_2018,filing_cabinet_200]=True
    inside[shampoo_2019,home_office_241]=True
    inside[pencil_2020,home_office_241]=True
    inside[food_food_2021,dining_room_41]=True
    inside[stamp_2022,home_office_241]=True
    inside[tea_bag_2023,bedroom_162]=True
    inside[ice_2024,dining_room_41]=True
    inside[ice_2024,sink_120]=True
    inside[rag_2025,bedroom_162]=True
    inside[rag_2025,filing_cabinet_200]=True
    inside[check_2026,bedroom_162]=True
    inside[food_orange_2027,dining_room_41]=True
    inside[instrument_guitar_2028,bedroom_162]=True
    inside[phone_2029,bathroom_1]=True
    inside[cd_2030,bedroom_162]=True
    inside[cd_2030,filing_cabinet_200]=True
    inside[scrabble_2031,bedroom_162]=True
    inside[scrabble_2031,filing_cabinet_200]=True
    inside[shoes_2033,home_office_241]=True
    inside[laser_pointer_2034,bedroom_162]=True
    inside[knife_2035,dining_room_41]=True
    inside[clothes_pants_2036,home_office_241]=True
    inside[knife_2037,dining_room_41]=True
    inside[knife_2037,cupboard_118]=True
    inside[box_2038,dining_room_41]=True
    inside[lighter_2039,dining_room_41]=True
    inside[pot_2040,dining_room_41]=True
    inside[pot_2040,microwave_135]=True
    inside[food_salt_2041,dining_room_41]=True
    inside[after_shave_2042,bedroom_162]=True
    inside[after_shave_2042,filing_cabinet_200]=True
    inside[stamp_2043,home_office_241]=True
    inside[shoe_rack_2044,bedroom_162]=True
    inside[glue_2045,dining_room_41]=True
    inside[glue_2045,trashcan_99]=True
    inside[food_food_2046,dining_room_41]=True
    inside[food_food_2046,fridge_126]=True
    inside[homework_2047,bedroom_162]=True
    inside[homework_2047,filing_cabinet_200]=True
    inside[food_onion_2048,dining_room_41]=True
    inside[food_onion_2048,fridge_126]=True
    inside[cup_2049,dining_room_41]=True
    inside[stereo_2050,bedroom_162]=True
    inside[stereo_2050,filing_cabinet_200]=True
    inside[after_shave_2051,bedroom_162]=True
    inside[after_shave_2051,filing_cabinet_200]=True
    inside[rag_2052,bedroom_162]=True
    inside[coffee_filter_2053,dining_room_41]=True
    inside[coffee_filter_2053,cupboard_117]=True
    inside[food_kiwi_2054,dining_room_41]=True
    inside[envelope_2055,dining_room_41]=True
    inside[toy_2056,bathroom_1]=True
    inside[blow_dryer_2057,home_office_241]=True
    inside[blow_dryer_2057,dresser_274]=True
    inside[check_2058,dining_room_41]=True
    inside[tooth_paste_2059,bathroom_1]=True
    inside[tooth_paste_2059,bathroom_cabinet_17]=True
    inside[novel_2060,bedroom_162]=True
    inside[food_orange_2061,dining_room_41]=True
    inside[food_orange_2061,trashcan_99]=True
    inside[piano_bench_2062,dining_room_41]=True
    inside[after_shave_2063,bathroom_1]=True
    inside[after_shave_2063,sink_19]=True
    inside[food_food_2064,dining_room_41]=True
    inside[coffee_filter_2065,dining_room_41]=True
    inside[coffee_filter_2065,coffe_maker_130]=True
    inside[tea_2066,dining_room_41]=True
    inside[tea_2066,cupboard_118]=True
    inside[piano_bench_2067,bathroom_1]=True
    inside[tray_2068,dining_room_41]=True
    inside[cat_2069,home_office_241]=True
    inside[cat_2069,dresser_274]=True
    inside[chessboard_2070,bedroom_162]=True
    inside[check_2071,bedroom_162]=True
    inside[food_cheese_2072,dining_room_41]=True
    inside[food_cheese_2072,oven_127]=True
    inside[food_food_2073,dining_room_41]=True
    inside[food_food_2073,fridge_126]=True
    inside[food_food_2074,bedroom_162]=True
    inside[food_food_2074,filing_cabinet_200]=True
    inside[check_2075,home_office_241]=True
    inside[check_2075,dresser_274]=True
    inside[toilet_paper_2076,bathroom_1]=True
    inside[toilet_paper_2076,toilet_15]=True
    inside[food_peanut_butter_2077,dining_room_41]=True
    inside[food_peanut_butter_2077,cupboard_118]=True
    between[door_38,bathroom_1]=True
    between[door_38,dining_room_41]=True
    between[door_61,dining_room_41]=True
    between[door_61,bedroom_162]=True
    between[door_62,dining_room_41]=True
    between[door_62,home_office_241]=True
    close[clothes_pants_2157,basket_for_clothes_2078]=True
    close[clothes_shirt_2158,basket_for_clothes_2078]=True
    close[clothes_socks_2159,basket_for_clothes_2078]=True
    close[clothes_skirt_2160,basket_for_clothes_2078]=True
    close[iron_2161,bowl_2142]=True
    close[basket_for_clothes_2078,clothes_pants_2157]=True
    close[basket_for_clothes_2078,clothes_shirt_2158]=True
    close[basket_for_clothes_2078,clothes_socks_2159]=True
    close[basket_for_clothes_2078,clothes_skirt_2160]=True
    close[basket_for_clothes_2078,sink_120]=True
    close[basket_for_clothes_2078,fridge_126]=True
    close[washing_machine_2079,sink_120]=True
    close[washing_machine_2079,fridge_126]=True
    close[food_steak_2080,fridge_126]=True
    close[food_apple_2081,fridge_126]=True
    close[food_bacon_2082,fridge_126]=True
    close[food_banana_2083,fridge_126]=True
    close[food_bread_2084,table_114]=True
    close[food_cake_2085,fridge_126]=True
    close[food_carrot_2086,fridge_126]=True
    close[food_cereal_2087,fridge_126]=True
    close[food_cheese_2088,fridge_126]=True
    close[food_chicken_2089,fridge_126]=True
    close[food_dessert_2090,fridge_126]=True
    close[food_donut_2091,fridge_126]=True
    close[food_egg_2092,fridge_126]=True
    close[food_fish_2093,fridge_126]=True
    close[food_food_2094,fridge_126]=True
    close[food_fruit_2095,fridge_126]=True
    close[food_hamburger_2096,fridge_126]=True
    close[food_ice_cream_2097,fridge_126]=True
    close[food_jam_2098,fridge_126]=True
    close[food_kiwi_2099,fridge_126]=True
    close[food_lemon_2100,fridge_126]=True
    close[food_noodles_2101,fridge_126]=True
    close[food_oatmeal_2102,fridge_126]=True
    close[food_orange_2103,fridge_126]=True
    close[food_onion_2104,fridge_126]=True
    close[food_peanut_butter_2105,fridge_126]=True
    close[food_pizza_2106,fridge_126]=True
    close[food_potato_2107,fridge_126]=True
    close[food_rice_2108,fridge_126]=True
    close[food_salt_2109,fridge_126]=True
    close[food_snack_2110,fridge_126]=True
    close[food_sugar_2111,fridge_126]=True
    close[food_turkey_2112,fridge_126]=True
    close[food_vegetable_2113,fridge_126]=True
    close[dry_pasta_2114,table_114]=True
    close[milk_2115,table_114]=True
    close[clothes_dress_2116,bed_197]=True
    close[clothes_hat_2117,table_114]=True
    close[clothes_gloves_2118,table_114]=True
    close[clothes_jacket_2119,couch_198]=True
    close[clothes_scarf_2120,bed_197]=True
    close[clothes_underwear_2121,bed_197]=True
    close[knife_2122,table_114]=True
    close[cutting_board_2123,kitchen_counter_119]=True
    close[remote_control_2124,tvstand_273]=True
    close[soap_2125,sink_19]=True
    close[soap_2126,sink_120]=True
    close[towel_2128,drawing_33]=True
    close[cd_player_2129,tvstand_273]=True
    close[dvd_player_2130,tvstand_273]=True
    close[headset_2131,tvstand_273]=True
    close[cup_2132,table_114]=True
    close[cup_2133,table_114]=True
    close[cup_2134,table_114]=True
    close[stove_2135,kitchen_counter_119]=True
    close[book_2136,bookshelf_124]=True
    close[book_2137,bookshelf_124]=True
    close[pot_2138,kitchen_counter_119]=True
    close[vacuum_cleaner_2139,trashcan_99]=True
    close[bowl_2140,kitchen_counter_119]=True
    close[bowl_2141,kitchen_counter_119]=True
    close[bowl_2142,iron_2161]=True
    close[bowl_2142,kitchen_counter_119]=True
    close[cleaning_solution_2143,sink_19]=True
    close[ironing_board_2144,dining_room_41]=True
    close[cd_2145,tvstand_273]=True
    close[headset_2146,desk_272]=True
    close[phone_2147,desk_272]=True
    close[sauce_2148,fridge_126]=True
    close[oil_2149,kitchen_counter_123]=True
    close[fork_2150,kitchen_counter_119]=True
    close[fork_2151,kitchen_counter_119]=True
    close[plate_2152,kitchen_counter_119]=True
    close[spectacles_2153,kitchen_counter_122]=True
    close[fryingpan_2154,kitchen_counter_122]=True
    close[detergent_2155,sink_19]=True
    close[window_2156,bathroom_1]=True
    close[bathroom_1,window_2156]=True
    close[wall_2,wall_3]=True
    close[wall_2,wall_5]=True
    close[wall_2,ceiling_6]=True
    close[wall_2,ceiling_7]=True
    close[wall_2,ceiling_8]=True
    close[wall_2,floor_10]=True
    close[wall_2,floor_11]=True
    close[wall_2,floor_12]=True
    close[wall_2,floor_13]=True
    close[wall_2,toilet_15]=True
    close[wall_2,shower_16]=True
    close[wall_2,curtain_22]=True
    close[wall_2,mat_32]=True
    close[wall_2,ceilinglamp_35]=True
    close[wall_2,doorjamb_37]=True
    close[wall_2,door_38]=True
    close[wall_2,light_39]=True
    close[wall_2,floor_42]=True
    close[wall_2,floor_43]=True
    close[wall_2,ceiling_52]=True
    close[wall_2,wall_63]=True
    close[wall_2,wall_70]=True
    close[wall_2,pillow_108]=True
    close[wall_2,drawing_111]=True
    close[wall_2,tvstand_116]=True
    close[wall_2,photoframe_219]=True
    close[wall_3,wall_2]=True
    close[wall_3,wall_4]=True
    close[wall_3,ceiling_6]=True
    close[wall_3,ceiling_7]=True
    close[wall_3,ceiling_9]=True
    close[wall_3,floor_10]=True
    close[wall_3,floor_11]=True
    close[wall_3,floor_12]=True
    close[wall_3,floor_14]=True
    close[wall_3,bathroom_cabinet_17]=True
    close[wall_3,bathroom_counter_18]=True
    close[wall_3,sink_19]=True
    close[wall_3,faucet_20]=True
    close[wall_3,mat_32]=True
    close[wall_3,walllamp_34]=True
    close[wall_3,ceilinglamp_35]=True
    close[wall_4,wall_3]=True
    close[wall_4,wall_5]=True
    close[wall_4,ceiling_6]=True
    close[wall_4,ceiling_8]=True
    close[wall_4,ceiling_9]=True
    close[wall_4,floor_10]=True
    close[wall_4,floor_11]=True
    close[wall_4,floor_13]=True
    close[wall_4,floor_14]=True
    close[wall_4,bathroom_cabinet_17]=True
    close[wall_4,bathroom_counter_18]=True
    close[wall_4,sink_19]=True
    close[wall_4,faucet_20]=True
    close[wall_4,curtain_22]=True
    close[wall_4,mat_32]=True
    close[wall_4,drawing_33]=True
    close[wall_4,ceilinglamp_35]=True
    close[wall_4,walllamp_36]=True
    close[wall_5,wall_2]=True
    close[wall_5,wall_4]=True
    close[wall_5,ceiling_7]=True
    close[wall_5,ceiling_8]=True
    close[wall_5,ceiling_9]=True
    close[wall_5,floor_12]=True
    close[wall_5,floor_13]=True
    close[wall_5,floor_14]=True
    close[wall_5,toilet_15]=True
    close[wall_5,shower_16]=True
    close[wall_5,shower_21]=True
    close[wall_5,curtain_22]=True
    close[wall_5,mat_32]=True
    close[wall_5,drawing_33]=True
    close[wall_5,ceilinglamp_35]=True
    close[wall_5,doorjamb_37]=True
    close[wall_5,door_38]=True
    close[wall_5,floor_170]=True
    close[wall_5,wall_174]=True
    close[wall_5,wall_176]=True
    close[wall_5,ceiling_183]=True
    close[wall_5,filing_cabinet_200]=True
    close[wall_5,drawing_202]=True
    close[wall_5,photoframe_219]=True
    close[ceiling_6,wall_2]=True
    close[ceiling_6,wall_3]=True
    close[ceiling_6,wall_4]=True
    close[ceiling_6,ceiling_7]=True
    close[ceiling_6,ceiling_9]=True
    close[ceiling_6,bathroom_cabinet_17]=True
    close[ceiling_6,faucet_20]=True
    close[ceiling_6,walllamp_34]=True
    close[ceiling_6,ceilinglamp_35]=True
    close[ceiling_7,wall_2]=True
    close[ceiling_7,wall_3]=True
    close[ceiling_7,wall_5]=True
    close[ceiling_7,ceiling_6]=True
    close[ceiling_7,ceiling_8]=True
    close[ceiling_7,shower_16]=True
    close[ceiling_7,ceilinglamp_35]=True
    close[ceiling_7,doorjamb_37]=True
    close[ceiling_7,light_39]=True
    close[ceiling_7,ceiling_52]=True
    close[ceiling_7,wall_70]=True
    close[ceiling_8,wall_2]=True
    close[ceiling_8,wall_4]=True
    close[ceiling_8,wall_5]=True
    close[ceiling_8,ceiling_7]=True
    close[ceiling_8,ceiling_9]=True
    close[ceiling_8,shower_16]=True
    close[ceiling_8,shower_21]=True
    close[ceiling_8,curtain_22]=True
    close[ceiling_8,drawing_33]=True
    close[ceiling_8,ceilinglamp_35]=True
    close[ceiling_8,wall_176]=True
    close[ceiling_8,ceiling_183]=True
    close[ceiling_8,drawing_202]=True
    close[ceiling_9,wall_3]=True
    close[ceiling_9,wall_4]=True
    close[ceiling_9,wall_5]=True
    close[ceiling_9,ceiling_6]=True
    close[ceiling_9,ceiling_8]=True
    close[ceiling_9,bathroom_cabinet_17]=True
    close[ceiling_9,faucet_20]=True
    close[ceiling_9,drawing_33]=True
    close[ceiling_9,ceilinglamp_35]=True
    close[ceiling_9,walllamp_36]=True
    close[floor_10,wall_2]=True
    close[floor_10,wall_3]=True
    close[floor_10,wall_4]=True
    close[floor_10,floor_11]=True
    close[floor_10,floor_12]=True
    close[floor_10,floor_14]=True
    close[floor_10,bathroom_counter_18]=True
    close[floor_10,sink_19]=True
    close[floor_10,faucet_20]=True
    close[floor_10,mat_32]=True
    close[floor_10,walllamp_34]=True
    close[floor_11,wall_2]=True
    close[floor_11,wall_3]=True
    close[floor_11,wall_4]=True
    close[floor_11,floor_10]=True
    close[floor_11,floor_12]=True
    close[floor_11,floor_14]=True
    close[floor_11,bathroom_counter_18]=True
    close[floor_11,sink_19]=True
    close[floor_11,faucet_20]=True
    close[floor_11,mat_32]=True
    close[floor_11,walllamp_34]=True
    close[floor_12,wall_2]=True
    close[floor_12,wall_3]=True
    close[floor_12,wall_5]=True
    close[floor_12,floor_10]=True
    close[floor_12,floor_11]=True
    close[floor_12,floor_13]=True
    close[floor_12,toilet_15]=True
    close[floor_12,shower_16]=True
    close[floor_12,mat_32]=True
    close[floor_12,doorjamb_37]=True
    close[floor_12,door_38]=True
    close[floor_12,light_39]=True
    close[floor_12,floor_42]=True
    close[floor_12,floor_43]=True
    close[floor_12,wall_70]=True
    close[floor_12,pillow_108]=True
    close[floor_12,tvstand_116]=True
    close[floor_12,photoframe_219]=True
    close[floor_13,wall_2]=True
    close[floor_13,wall_4]=True
    close[floor_13,wall_5]=True
    close[floor_13,floor_12]=True
    close[floor_13,floor_14]=True
    close[floor_13,toilet_15]=True
    close[floor_13,shower_16]=True
    close[floor_13,shower_21]=True
    close[floor_13,curtain_22]=True
    close[floor_13,mat_32]=True
    close[floor_13,door_38]=True
    close[floor_13,floor_170]=True
    close[floor_13,wall_176]=True
    close[floor_13,filing_cabinet_200]=True
    close[floor_13,photoframe_219]=True
    close[floor_14,wall_3]=True
    close[floor_14,wall_4]=True
    close[floor_14,wall_5]=True
    close[floor_14,floor_10]=True
    close[floor_14,floor_11]=True
    close[floor_14,floor_13]=True
    close[floor_14,bathroom_counter_18]=True
    close[floor_14,sink_19]=True
    close[floor_14,faucet_20]=True
    close[floor_14,mat_32]=True
    close[floor_14,drawing_33]=True
    close[floor_14,walllamp_36]=True
    close[toilet_15,wall_2]=True
    close[toilet_15,wall_5]=True
    close[toilet_15,floor_12]=True
    close[toilet_15,floor_13]=True
    close[toilet_15,shower_16]=True
    close[toilet_15,shower_21]=True
    close[toilet_15,curtain_22]=True
    close[toilet_15,doorjamb_37]=True
    close[toilet_15,door_38]=True
    close[toilet_15,floor_42]=True
    close[toilet_15,floor_43]=True
    close[toilet_15,wall_70]=True
    close[toilet_15,floor_170]=True
    close[toilet_15,wall_176]=True
    close[toilet_15,bookshelf_196]=True
    close[toilet_15,filing_cabinet_200]=True
    close[toilet_15,photoframe_219]=True
    close[toilet_15,toilet_paper_2076]=True
    close[shower_16,wall_2]=True
    close[shower_16,wall_5]=True
    close[shower_16,ceiling_7]=True
    close[shower_16,ceiling_8]=True
    close[shower_16,floor_12]=True
    close[shower_16,floor_13]=True
    close[shower_16,toilet_15]=True
    close[shower_16,shower_21]=True
    close[shower_16,curtain_22]=True
    close[shower_16,mat_32]=True
    close[shower_16,ceilinglamp_35]=True
    close[shower_16,doorjamb_37]=True
    close[shower_16,door_38]=True
    close[shower_16,light_39]=True
    close[shower_16,floor_42]=True
    close[shower_16,floor_43]=True
    close[shower_16,ceiling_52]=True
    close[shower_16,wall_70]=True
    close[shower_16,floor_170]=True
    close[shower_16,wall_176]=True
    close[shower_16,ceiling_183]=True
    close[shower_16,bookshelf_196]=True
    close[shower_16,filing_cabinet_200]=True
    close[shower_16,photoframe_219]=True
    close[bathroom_cabinet_17,wall_3]=True
    close[bathroom_cabinet_17,wall_4]=True
    close[bathroom_cabinet_17,ceiling_6]=True
    close[bathroom_cabinet_17,ceiling_9]=True
    close[bathroom_cabinet_17,bathroom_counter_18]=True
    close[bathroom_cabinet_17,sink_19]=True
    close[bathroom_cabinet_17,faucet_20]=True
    close[bathroom_cabinet_17,walllamp_34]=True
    close[bathroom_cabinet_17,walllamp_36]=True
    close[bathroom_cabinet_17,tooth_paste_2059]=True
    close[bathroom_counter_18,wall_3]=True
    close[bathroom_counter_18,wall_4]=True
    close[bathroom_counter_18,floor_10]=True
    close[bathroom_counter_18,floor_11]=True
    close[bathroom_counter_18,floor_14]=True
    close[bathroom_counter_18,bathroom_cabinet_17]=True
    close[bathroom_counter_18,sink_19]=True
    close[bathroom_counter_18,faucet_20]=True
    close[bathroom_counter_18,mat_32]=True
    close[bathroom_counter_18,walllamp_34]=True
    close[bathroom_counter_18,walllamp_36]=True
    close[bathroom_counter_18,phone_2029]=True
    close[sink_19,soap_2125]=True
    close[sink_19,cleaning_solution_2143]=True
    close[sink_19,detergent_2155]=True
    close[sink_19,wall_3]=True
    close[sink_19,wall_4]=True
    close[sink_19,floor_10]=True
    close[sink_19,floor_11]=True
    close[sink_19,floor_14]=True
    close[sink_19,bathroom_cabinet_17]=True
    close[sink_19,bathroom_counter_18]=True
    close[sink_19,faucet_20]=True
    close[sink_19,mat_32]=True
    close[sink_19,after_shave_2063]=True
    close[faucet_20,wall_3]=True
    close[faucet_20,wall_4]=True
    close[faucet_20,ceiling_6]=True
    close[faucet_20,ceiling_9]=True
    close[faucet_20,floor_10]=True
    close[faucet_20,floor_11]=True
    close[faucet_20,floor_14]=True
    close[faucet_20,bathroom_cabinet_17]=True
    close[faucet_20,bathroom_counter_18]=True
    close[faucet_20,sink_19]=True
    close[faucet_20,mat_32]=True
    close[shower_21,wall_5]=True
    close[shower_21,ceiling_8]=True
    close[shower_21,floor_13]=True
    close[shower_21,toilet_15]=True
    close[shower_21,shower_16]=True
    close[shower_21,curtain_22]=True
    close[shower_21,ceilinglamp_35]=True
    close[shower_21,floor_170]=True
    close[shower_21,wall_174]=True
    close[shower_21,wall_176]=True
    close[shower_21,ceiling_183]=True
    close[shower_21,filing_cabinet_200]=True
    close[shower_21,drawing_202]=True
    close[shower_21,photoframe_219]=True
    close[curtain_22,wall_2]=True
    close[curtain_22,wall_4]=True
    close[curtain_22,wall_5]=True
    close[curtain_22,ceiling_8]=True
    close[curtain_22,floor_13]=True
    close[curtain_22,toilet_15]=True
    close[curtain_22,shower_16]=True
    close[curtain_22,shower_21]=True
    close[curtain_22,mat_32]=True
    close[curtain_22,ceilinglamp_35]=True
    close[mat_32,wall_2]=True
    close[mat_32,wall_3]=True
    close[mat_32,wall_4]=True
    close[mat_32,wall_5]=True
    close[mat_32,floor_10]=True
    close[mat_32,floor_11]=True
    close[mat_32,floor_12]=True
    close[mat_32,floor_13]=True
    close[mat_32,floor_14]=True
    close[mat_32,shower_16]=True
    close[mat_32,bathroom_counter_18]=True
    close[mat_32,sink_19]=True
    close[mat_32,faucet_20]=True
    close[mat_32,curtain_22]=True
    close[mat_32,toy_2056]=True
    close[mat_32,piano_bench_2067]=True
    close[drawing_33,towel_2128]=True
    close[drawing_33,wall_4]=True
    close[drawing_33,wall_5]=True
    close[drawing_33,ceiling_8]=True
    close[drawing_33,ceiling_9]=True
    close[drawing_33,floor_14]=True
    close[drawing_33,walllamp_36]=True
    close[walllamp_34,wall_3]=True
    close[walllamp_34,ceiling_6]=True
    close[walllamp_34,floor_10]=True
    close[walllamp_34,floor_11]=True
    close[walllamp_34,bathroom_cabinet_17]=True
    close[walllamp_34,bathroom_counter_18]=True
    close[ceilinglamp_35,wall_2]=True
    close[ceilinglamp_35,wall_3]=True
    close[ceilinglamp_35,wall_4]=True
    close[ceilinglamp_35,wall_5]=True
    close[ceilinglamp_35,ceiling_6]=True
    close[ceilinglamp_35,ceiling_7]=True
    close[ceilinglamp_35,ceiling_8]=True
    close[ceilinglamp_35,ceiling_9]=True
    close[ceilinglamp_35,shower_16]=True
    close[ceilinglamp_35,shower_21]=True
    close[ceilinglamp_35,curtain_22]=True
    close[walllamp_36,wall_4]=True
    close[walllamp_36,ceiling_9]=True
    close[walllamp_36,floor_14]=True
    close[walllamp_36,bathroom_cabinet_17]=True
    close[walllamp_36,bathroom_counter_18]=True
    close[walllamp_36,drawing_33]=True
    close[doorjamb_37,wall_2]=True
    close[doorjamb_37,wall_5]=True
    close[doorjamb_37,ceiling_7]=True
    close[doorjamb_37,floor_12]=True
    close[doorjamb_37,toilet_15]=True
    close[doorjamb_37,shower_16]=True
    close[doorjamb_37,door_38]=True
    close[doorjamb_37,light_39]=True
    close[doorjamb_37,floor_42]=True
    close[doorjamb_37,floor_43]=True
    close[doorjamb_37,ceiling_52]=True
    close[doorjamb_37,wall_63]=True
    close[doorjamb_37,wall_70]=True
    close[doorjamb_37,pillow_108]=True
    close[doorjamb_37,bookshelf_124]=True
    close[doorjamb_37,wall_176]=True
    close[doorjamb_37,bookshelf_196]=True
    close[doorjamb_37,photoframe_219]=True
    close[door_38,wall_2]=True
    close[door_38,wall_5]=True
    close[door_38,floor_12]=True
    close[door_38,floor_13]=True
    close[door_38,toilet_15]=True
    close[door_38,shower_16]=True
    close[door_38,doorjamb_37]=True
    close[door_38,light_39]=True
    close[door_38,floor_42]=True
    close[door_38,floor_43]=True
    close[door_38,floor_48]=True
    close[door_38,wall_63]=True
    close[door_38,wall_70]=True
    close[door_38,pillow_108]=True
    close[door_38,drawing_110]=True
    close[door_38,tvstand_116]=True
    close[door_38,bookshelf_124]=True
    close[door_38,floor_170]=True
    close[door_38,wall_176]=True
    close[door_38,bookshelf_196]=True
    close[door_38,photoframe_219]=True
    close[light_39,wall_2]=True
    close[light_39,ceiling_7]=True
    close[light_39,floor_12]=True
    close[light_39,shower_16]=True
    close[light_39,doorjamb_37]=True
    close[light_39,door_38]=True
    close[light_39,floor_42]=True
    close[light_39,floor_43]=True
    close[light_39,floor_48]=True
    close[light_39,ceiling_52]=True
    close[light_39,ceiling_57]=True
    close[light_39,wall_63]=True
    close[light_39,wall_70]=True
    close[light_39,pillow_108]=True
    close[light_39,drawing_111]=True
    close[light_39,tvstand_116]=True
    close[dining_room_41,ironing_board_2144]=True
    close[floor_42,wall_2]=True
    close[floor_42,floor_12]=True
    close[floor_42,toilet_15]=True
    close[floor_42,shower_16]=True
    close[floor_42,doorjamb_37]=True
    close[floor_42,door_38]=True
    close[floor_42,light_39]=True
    close[floor_42,floor_43]=True
    close[floor_42,floor_44]=True
    close[floor_42,floor_48]=True
    close[floor_42,door_61]=True
    close[floor_42,wall_70]=True
    close[floor_42,powersocket_72]=True
    close[floor_42,mat_102]=True
    close[floor_42,pillow_106]=True
    close[floor_42,pillow_108]=True
    close[floor_42,bench_115]=True
    close[floor_42,tvstand_116]=True
    close[floor_42,bookshelf_124]=True
    close[floor_42,floor_170]=True
    close[floor_42,wall_176]=True
    close[floor_42,bookshelf_196]=True
    close[floor_42,light_212]=True
    close[floor_42,photoframe_219]=True
    close[floor_43,wall_2]=True
    close[floor_43,floor_12]=True
    close[floor_43,toilet_15]=True
    close[floor_43,shower_16]=True
    close[floor_43,doorjamb_37]=True
    close[floor_43,door_38]=True
    close[floor_43,light_39]=True
    close[floor_43,floor_42]=True
    close[floor_43,floor_44]=True
    close[floor_43,floor_48]=True
    close[floor_43,door_61]=True
    close[floor_43,wall_70]=True
    close[floor_43,powersocket_72]=True
    close[floor_43,mat_102]=True
    close[floor_43,pillow_106]=True
    close[floor_43,pillow_108]=True
    close[floor_43,bench_115]=True
    close[floor_43,tvstand_116]=True
    close[floor_43,bookshelf_124]=True
    close[floor_43,floor_170]=True
    close[floor_43,wall_176]=True
    close[floor_43,bookshelf_196]=True
    close[floor_43,light_212]=True
    close[floor_43,photoframe_219]=True
    close[floor_44,floor_42]=True
    close[floor_44,floor_43]=True
    close[floor_44,floor_45]=True
    close[floor_44,floor_47]=True
    close[floor_44,door_61]=True
    close[floor_44,wall_66]=True
    close[floor_44,wall_67]=True
    close[floor_44,wall_70]=True
    close[floor_44,powersocket_72]=True
    close[floor_44,light_73]=True
    close[floor_44,mat_102]=True
    close[floor_44,pillow_104]=True
    close[floor_44,pillow_106]=True
    close[floor_44,bench_113]=True
    close[floor_44,table_114]=True
    close[floor_44,bench_115]=True
    close[floor_44,bookshelf_124]=True
    close[floor_44,fridge_126]=True
    close[floor_44,floor_169]=True
    close[floor_44,wall_179]=True
    close[floor_44,doorjamb_190]=True
    close[floor_44,desk_193]=True
    close[floor_44,bookshelf_196]=True
    close[floor_44,computer_209]=True
    close[floor_44,light_212]=True
    close[floor_44,mouse_213]=True
    close[floor_44,mousepad_214]=True
    close[floor_44,piano_bench_2006]=True
    close[floor_44,piano_bench_2062]=True
    close[floor_45,floor_44]=True
    close[floor_45,floor_46]=True
    close[floor_45,door_61]=True
    close[floor_45,wall_67]=True
    close[floor_45,light_73]=True
    close[floor_45,knifeblock_76]=True
    close[floor_45,pillow_104]=True
    close[floor_45,bench_113]=True
    close[floor_45,kitchen_counter_119]=True
    close[floor_45,sink_120]=True
    close[floor_45,faucet_121]=True
    close[floor_45,kitchen_counter_123]=True
    close[floor_45,fridge_126]=True
    close[floor_45,floor_163]=True
    close[floor_45,floor_164]=True
    close[floor_45,wall_175]=True
    close[floor_45,desk_193]=True
    close[floor_45,computer_209]=True
    close[floor_45,cpuscreen_210]=True
    close[floor_45,keyboard_211]=True
    close[floor_45,mouse_213]=True
    close[floor_45,mousepad_214]=True
    close[floor_46,floor_45]=True
    close[floor_46,floor_47]=True
    close[floor_46,floor_51]=True
    close[floor_46,wall_64]=True
    close[floor_46,wall_67]=True
    close[floor_46,wall_68]=True
    close[floor_46,knifeblock_76]=True
    close[floor_46,pot_78]=True
    close[floor_46,mat_102]=True
    close[floor_46,pillow_103]=True
    close[floor_46,pillow_104]=True
    close[floor_46,bench_113]=True
    close[floor_46,kitchen_counter_119]=True
    close[floor_46,sink_120]=True
    close[floor_46,faucet_121]=True
    close[floor_46,kitchen_counter_122]=True
    close[floor_46,oven_127]=True
    close[floor_46,tray_128]=True
    close[floor_46,dishwasher_129]=True
    close[floor_46,toaster_132]=True
    close[floor_47,floor_44]=True
    close[floor_47,floor_46]=True
    close[floor_47,floor_48]=True
    close[floor_47,floor_50]=True
    close[floor_47,mat_102]=True
    close[floor_47,pillow_103]=True
    close[floor_47,pillow_104]=True
    close[floor_47,pillow_105]=True
    close[floor_47,pillow_106]=True
    close[floor_47,bench_113]=True
    close[floor_47,table_114]=True
    close[floor_47,bench_115]=True
    close[floor_48,door_38]=True
    close[floor_48,light_39]=True
    close[floor_48,floor_42]=True
    close[floor_48,floor_43]=True
    close[floor_48,floor_47]=True
    close[floor_48,floor_49]=True
    close[floor_48,wall_63]=True
    close[floor_48,wall_69]=True
    close[floor_48,wall_70]=True
    close[floor_48,mat_102]=True
    close[floor_48,pillow_105]=True
    close[floor_48,pillow_106]=True
    close[floor_48,pillow_107]=True
    close[floor_48,pillow_108]=True
    close[floor_48,drawing_111]=True
    close[floor_48,table_114]=True
    close[floor_48,bench_115]=True
    close[floor_48,tvstand_116]=True
    close[floor_49,floor_48]=True
    close[floor_49,floor_50]=True
    close[floor_49,door_62]=True
    close[floor_49,wall_69]=True
    close[floor_49,phone_71]=True
    close[floor_49,mat_102]=True
    close[floor_49,pillow_105]=True
    close[floor_49,pillow_107]=True
    close[floor_49,bench_115]=True
    close[floor_49,tvstand_116]=True
    close[floor_49,wall_244]=True
    close[floor_49,floor_261]=True
    close[floor_49,tvstand_273]=True
    close[floor_49,powersocket_282]=True
    close[floor_49,light_283]=True
    close[floor_49,mat_284]=True
    close[floor_49,doorjamb_309]=True
    close[floor_50,floor_47]=True
    close[floor_50,floor_49]=True
    close[floor_50,floor_51]=True
    close[floor_50,door_62]=True
    close[floor_50,wall_65]=True
    close[floor_50,wall_68]=True
    close[floor_50,wall_69]=True
    close[floor_50,trashcan_99]=True
    close[floor_50,mat_102]=True
    close[floor_50,pillow_103]=True
    close[floor_50,pillow_105]=True
    close[floor_50,bench_113]=True
    close[floor_50,table_114]=True
    close[floor_50,bench_115]=True
    close[floor_50,wall_246]=True
    close[floor_50,floor_262]=True
    close[floor_50,bookshelf_275]=True
    close[floor_50,light_283]=True
    close[floor_51,floor_46]=True
    close[floor_51,floor_50]=True
    close[floor_51,wall_68]=True
    close[floor_51,trashcan_99]=True
    close[floor_51,pillow_103]=True
    close[floor_51,bench_113]=True
    close[floor_51,kitchen_counter_122]=True
    close[floor_51,oven_127]=True
    close[floor_51,tray_128]=True
    close[floor_51,dishwasher_129]=True
    close[floor_51,coffe_maker_130]=True
    close[floor_51,toaster_132]=True
    close[floor_51,microwave_135]=True
    close[floor_51,bookshelf_275]=True
    close[ceiling_52,wall_2]=True
    close[ceiling_52,ceiling_7]=True
    close[ceiling_52,shower_16]=True
    close[ceiling_52,doorjamb_37]=True
    close[ceiling_52,light_39]=True
    close[ceiling_52,ceiling_53]=True
    close[ceiling_52,ceiling_57]=True
    close[ceiling_52,wall_70]=True
    close[ceiling_52,drawing_110]=True
    close[ceiling_52,ceilinglamp_137]=True
    close[ceiling_52,wall_176]=True
    close[ceiling_52,ceiling_183]=True
    close[ceiling_52,bookshelf_196]=True
    close[ceiling_52,light_212]=True
    close[ceiling_53,ceiling_52]=True
    close[ceiling_53,ceiling_54]=True
    close[ceiling_53,ceiling_56]=True
    close[ceiling_53,wall_66]=True
    close[ceiling_53,wall_67]=True
    close[ceiling_53,wall_70]=True
    close[ceiling_53,light_73]=True
    close[ceiling_53,drawing_110]=True
    close[ceiling_53,fridge_126]=True
    close[ceiling_53,ceilinglamp_137]=True
    close[ceiling_53,wall_179]=True
    close[ceiling_53,ceiling_182]=True
    close[ceiling_53,doorjamb_190]=True
    close[ceiling_53,light_212]=True
    close[ceiling_54,ceiling_53]=True
    close[ceiling_54,ceiling_55]=True
    close[ceiling_54,wall_67]=True
    close[ceiling_54,knifeblock_76]=True
    close[ceiling_54,cupboard_117]=True
    close[ceiling_54,faucet_121]=True
    close[ceiling_54,stovefan_125]=True
    close[ceiling_54,fridge_126]=True
    close[ceiling_54,ceilinglamp_137]=True
    close[ceiling_54,walllamp_140]=True
    close[ceiling_54,wall_175]=True
    close[ceiling_54,ceiling_181]=True
    close[ceiling_54,cpuscreen_210]=True
    close[ceiling_55,ceiling_54]=True
    close[ceiling_55,ceiling_56]=True
    close[ceiling_55,ceiling_60]=True
    close[ceiling_55,wall_64]=True
    close[ceiling_55,wall_67]=True
    close[ceiling_55,wall_68]=True
    close[ceiling_55,knifeblock_76]=True
    close[ceiling_55,pot_78]=True
    close[ceiling_55,cupboard_117]=True
    close[ceiling_55,cupboard_118]=True
    close[ceiling_55,stovefan_125]=True
    close[ceiling_55,oven_127]=True
    close[ceiling_55,toaster_132]=True
    close[ceiling_55,ceilinglamp_137]=True
    close[ceiling_55,ceilinglamp_138]=True
    close[ceiling_55,walllamp_139]=True
    close[ceiling_55,walllamp_140]=True
    close[ceiling_55,walllamp_141]=True
    close[ceiling_56,ceiling_53]=True
    close[ceiling_56,ceiling_55]=True
    close[ceiling_56,ceiling_57]=True
    close[ceiling_56,ceiling_59]=True
    close[ceiling_56,ceilinglamp_137]=True
    close[ceiling_56,ceilinglamp_138]=True
    close[ceiling_57,light_39]=True
    close[ceiling_57,ceiling_52]=True
    close[ceiling_57,ceiling_56]=True
    close[ceiling_57,ceiling_58]=True
    close[ceiling_57,wall_63]=True
    close[ceiling_57,wall_69]=True
    close[ceiling_57,wall_70]=True
    close[ceiling_57,phone_71]=True
    close[ceiling_57,drawing_111]=True
    close[ceiling_57,ceilinglamp_137]=True
    close[ceiling_57,ceilinglamp_138]=True
    close[ceiling_58,ceiling_57]=True
    close[ceiling_58,ceiling_59]=True
    close[ceiling_58,wall_69]=True
    close[ceiling_58,phone_71]=True
    close[ceiling_58,ceilinglamp_138]=True
    close[ceiling_58,wall_244]=True
    close[ceiling_58,ceiling_251]=True
    close[ceiling_58,light_283]=True
    close[ceiling_58,doorjamb_309]=True
    close[ceiling_59,ceiling_56]=True
    close[ceiling_59,ceiling_58]=True
    close[ceiling_59,ceiling_60]=True
    close[ceiling_59,wall_65]=True
    close[ceiling_59,wall_68]=True
    close[ceiling_59,wall_69]=True
    close[ceiling_59,ceilinglamp_138]=True
    close[ceiling_59,wall_246]=True
    close[ceiling_59,ceiling_252]=True
    close[ceiling_59,bookshelf_275]=True
    close[ceiling_60,ceiling_55]=True
    close[ceiling_60,ceiling_59]=True
    close[ceiling_60,wall_68]=True
    close[ceiling_60,cupboard_118]=True
    close[ceiling_60,stovefan_125]=True
    close[ceiling_60,coffe_maker_130]=True
    close[ceiling_60,toaster_132]=True
    close[ceiling_60,microwave_135]=True
    close[ceiling_60,ceilinglamp_138]=True
    close[ceiling_60,walllamp_139]=True
    close[ceiling_60,walllamp_141]=True
    close[door_61,floor_42]=True
    close[door_61,floor_43]=True
    close[door_61,floor_44]=True
    close[door_61,floor_45]=True
    close[door_61,wall_66]=True
    close[door_61,wall_67]=True
    close[door_61,wall_70]=True
    close[door_61,powersocket_72]=True
    close[door_61,light_73]=True
    close[door_61,fridge_126]=True
    close[door_61,floor_163]=True
    close[door_61,floor_164]=True
    close[door_61,floor_169]=True
    close[door_61,floor_170]=True
    close[door_61,wall_175]=True
    close[door_61,wall_176]=True
    close[door_61,wall_179]=True
    close[door_61,doorjamb_190]=True
    close[door_61,desk_193]=True
    close[door_61,bookshelf_196]=True
    close[door_61,computer_209]=True
    close[door_61,light_212]=True
    close[door_61,mouse_213]=True
    close[door_61,mousepad_214]=True
    close[door_62,floor_49]=True
    close[door_62,floor_50]=True
    close[door_62,wall_65]=True
    close[door_62,wall_69]=True
    close[door_62,phone_71]=True
    close[door_62,wall_244]=True
    close[door_62,wall_246]=True
    close[door_62,wall_247]=True
    close[door_62,floor_259]=True
    close[door_62,floor_260]=True
    close[door_62,floor_261]=True
    close[door_62,floor_262]=True
    close[door_62,tvstand_273]=True
    close[door_62,television_281]=True
    close[door_62,powersocket_282]=True
    close[door_62,light_283]=True
    close[door_62,mat_284]=True
    close[door_62,doorjamb_309]=True
    close[wall_63,wall_2]=True
    close[wall_63,doorjamb_37]=True
    close[wall_63,door_38]=True
    close[wall_63,light_39]=True
    close[wall_63,floor_48]=True
    close[wall_63,ceiling_57]=True
    close[wall_63,wall_69]=True
    close[wall_63,wall_70]=True
    close[wall_63,phone_71]=True
    close[wall_63,pillow_107]=True
    close[wall_63,pillow_108]=True
    close[wall_63,drawing_111]=True
    close[wall_63,tvstand_116]=True
    close[wall_64,floor_46]=True
    close[wall_64,ceiling_55]=True
    close[wall_64,wall_67]=True
    close[wall_64,wall_68]=True
    close[wall_64,knifeblock_76]=True
    close[wall_64,pot_78]=True
    close[wall_64,cupboard_117]=True
    close[wall_64,cupboard_118]=True
    close[wall_64,kitchen_counter_119]=True
    close[wall_64,sink_120]=True
    close[wall_64,faucet_121]=True
    close[wall_64,kitchen_counter_122]=True
    close[wall_64,stovefan_125]=True
    close[wall_64,oven_127]=True
    close[wall_64,tray_128]=True
    close[wall_64,dishwasher_129]=True
    close[wall_64,toaster_132]=True
    close[wall_64,microwave_135]=True
    close[wall_64,walllamp_139]=True
    close[wall_64,walllamp_140]=True
    close[wall_64,walllamp_141]=True
    close[wall_65,floor_50]=True
    close[wall_65,ceiling_59]=True
    close[wall_65,door_62]=True
    close[wall_65,wall_68]=True
    close[wall_65,wall_69]=True
    close[wall_65,trashcan_99]=True
    close[wall_65,wall_244]=True
    close[wall_65,wall_246]=True
    close[wall_65,ceiling_252]=True
    close[wall_65,floor_262]=True
    close[wall_65,bookshelf_275]=True
    close[wall_65,light_283]=True
    close[wall_65,doorjamb_309]=True
    close[wall_66,floor_44]=True
    close[wall_66,ceiling_53]=True
    close[wall_66,door_61]=True
    close[wall_66,wall_67]=True
    close[wall_66,wall_70]=True
    close[wall_66,powersocket_72]=True
    close[wall_66,light_73]=True
    close[wall_66,drawing_110]=True
    close[wall_66,bookshelf_124]=True
    close[wall_66,fridge_126]=True
    close[wall_66,floor_169]=True
    close[wall_66,wall_175]=True
    close[wall_66,wall_176]=True
    close[wall_66,wall_179]=True
    close[wall_66,ceiling_182]=True
    close[wall_66,doorjamb_190]=True
    close[wall_66,desk_193]=True
    close[wall_66,bookshelf_196]=True
    close[wall_66,computer_209]=True
    close[wall_66,cpuscreen_210]=True
    close[wall_66,keyboard_211]=True
    close[wall_66,light_212]=True
    close[wall_66,mouse_213]=True
    close[wall_66,mousepad_214]=True
    close[wall_67,floor_44]=True
    close[wall_67,floor_45]=True
    close[wall_67,floor_46]=True
    close[wall_67,ceiling_53]=True
    close[wall_67,ceiling_54]=True
    close[wall_67,ceiling_55]=True
    close[wall_67,door_61]=True
    close[wall_67,wall_64]=True
    close[wall_67,wall_66]=True
    close[wall_67,light_73]=True
    close[wall_67,knifeblock_76]=True
    close[wall_67,pot_78]=True
    close[wall_67,pillow_104]=True
    close[wall_67,bench_113]=True
    close[wall_67,cupboard_117]=True
    close[wall_67,kitchen_counter_119]=True
    close[wall_67,sink_120]=True
    close[wall_67,faucet_121]=True
    close[wall_67,kitchen_counter_123]=True
    close[wall_67,stovefan_125]=True
    close[wall_67,fridge_126]=True
    close[wall_67,oven_127]=True
    close[wall_67,tray_128]=True
    close[wall_67,ceilinglamp_137]=True
    close[wall_67,walllamp_140]=True
    close[wall_67,walllamp_141]=True
    close[wall_67,floor_163]=True
    close[wall_67,floor_164]=True
    close[wall_67,wall_175]=True
    close[wall_67,wall_179]=True
    close[wall_67,ceiling_181]=True
    close[wall_67,doorjamb_190]=True
    close[wall_67,desk_193]=True
    close[wall_67,computer_209]=True
    close[wall_67,cpuscreen_210]=True
    close[wall_67,keyboard_211]=True
    close[wall_67,mouse_213]=True
    close[wall_67,mousepad_214]=True
    close[wall_68,floor_46]=True
    close[wall_68,floor_50]=True
    close[wall_68,floor_51]=True
    close[wall_68,ceiling_55]=True
    close[wall_68,ceiling_59]=True
    close[wall_68,ceiling_60]=True
    close[wall_68,wall_64]=True
    close[wall_68,wall_65]=True
    close[wall_68,pot_78]=True
    close[wall_68,trashcan_99]=True
    close[wall_68,pillow_103]=True
    close[wall_68,bench_113]=True
    close[wall_68,cupboard_118]=True
    close[wall_68,kitchen_counter_122]=True
    close[wall_68,stovefan_125]=True
    close[wall_68,oven_127]=True
    close[wall_68,tray_128]=True
    close[wall_68,dishwasher_129]=True
    close[wall_68,coffe_maker_130]=True
    close[wall_68,toaster_132]=True
    close[wall_68,microwave_135]=True
    close[wall_68,ceilinglamp_138]=True
    close[wall_68,walllamp_139]=True
    close[wall_68,walllamp_141]=True
    close[wall_68,bookshelf_275]=True
    close[wall_69,floor_48]=True
    close[wall_69,floor_49]=True
    close[wall_69,floor_50]=True
    close[wall_69,ceiling_57]=True
    close[wall_69,ceiling_58]=True
    close[wall_69,ceiling_59]=True
    close[wall_69,door_62]=True
    close[wall_69,wall_63]=True
    close[wall_69,wall_65]=True
    close[wall_69,phone_71]=True
    close[wall_69,pillow_105]=True
    close[wall_69,pillow_107]=True
    close[wall_69,drawing_111]=True
    close[wall_69,bench_115]=True
    close[wall_69,tvstand_116]=True
    close[wall_69,ceilinglamp_138]=True
    close[wall_69,wall_244]=True
    close[wall_69,ceiling_251]=True
    close[wall_69,floor_261]=True
    close[wall_69,tvstand_273]=True
    close[wall_69,television_281]=True
    close[wall_69,powersocket_282]=True
    close[wall_69,light_283]=True
    close[wall_69,mat_284]=True
    close[wall_69,doorjamb_309]=True
    close[wall_70,wall_2]=True
    close[wall_70,ceiling_7]=True
    close[wall_70,floor_12]=True
    close[wall_70,toilet_15]=True
    close[wall_70,shower_16]=True
    close[wall_70,doorjamb_37]=True
    close[wall_70,door_38]=True
    close[wall_70,light_39]=True
    close[wall_70,floor_42]=True
    close[wall_70,floor_43]=True
    close[wall_70,floor_44]=True
    close[wall_70,floor_48]=True
    close[wall_70,ceiling_52]=True
    close[wall_70,ceiling_53]=True
    close[wall_70,ceiling_57]=True
    close[wall_70,door_61]=True
    close[wall_70,wall_63]=True
    close[wall_70,wall_66]=True
    close[wall_70,powersocket_72]=True
    close[wall_70,pillow_106]=True
    close[wall_70,pillow_108]=True
    close[wall_70,drawing_110]=True
    close[wall_70,drawing_111]=True
    close[wall_70,bench_115]=True
    close[wall_70,tvstand_116]=True
    close[wall_70,bookshelf_124]=True
    close[wall_70,ceilinglamp_137]=True
    close[wall_70,floor_170]=True
    close[wall_70,wall_176]=True
    close[wall_70,wall_179]=True
    close[wall_70,ceiling_183]=True
    close[wall_70,doorjamb_190]=True
    close[wall_70,bookshelf_196]=True
    close[wall_70,filing_cabinet_200]=True
    close[wall_70,light_212]=True
    close[wall_70,photoframe_219]=True
    close[phone_71,floor_49]=True
    close[phone_71,ceiling_57]=True
    close[phone_71,ceiling_58]=True
    close[phone_71,door_62]=True
    close[phone_71,wall_63]=True
    close[phone_71,wall_69]=True
    close[phone_71,pillow_107]=True
    close[phone_71,drawing_111]=True
    close[phone_71,tvstand_116]=True
    close[powersocket_72,floor_42]=True
    close[powersocket_72,floor_43]=True
    close[powersocket_72,floor_44]=True
    close[powersocket_72,door_61]=True
    close[powersocket_72,wall_66]=True
    close[powersocket_72,wall_70]=True
    close[powersocket_72,light_73]=True
    close[powersocket_72,bookshelf_124]=True
    close[powersocket_72,fridge_126]=True
    close[powersocket_72,floor_169]=True
    close[powersocket_72,floor_170]=True
    close[powersocket_72,wall_176]=True
    close[powersocket_72,wall_179]=True
    close[powersocket_72,doorjamb_190]=True
    close[powersocket_72,bookshelf_196]=True
    close[powersocket_72,light_212]=True
    close[light_73,floor_44]=True
    close[light_73,floor_45]=True
    close[light_73,ceiling_53]=True
    close[light_73,door_61]=True
    close[light_73,wall_66]=True
    close[light_73,wall_67]=True
    close[light_73,powersocket_72]=True
    close[light_73,fridge_126]=True
    close[light_73,floor_163]=True
    close[light_73,floor_164]=True
    close[light_73,floor_169]=True
    close[light_73,wall_175]=True
    close[light_73,wall_179]=True
    close[light_73,ceiling_182]=True
    close[light_73,doorjamb_190]=True
    close[light_73,desk_193]=True
    close[light_73,computer_209]=True
    close[light_73,cpuscreen_210]=True
    close[light_73,keyboard_211]=True
    close[light_73,light_212]=True
    close[light_73,mouse_213]=True
    close[light_73,mousepad_214]=True
    close[knifeblock_76,floor_45]=True
    close[knifeblock_76,floor_46]=True
    close[knifeblock_76,ceiling_54]=True
    close[knifeblock_76,ceiling_55]=True
    close[knifeblock_76,wall_64]=True
    close[knifeblock_76,wall_67]=True
    close[knifeblock_76,pot_78]=True
    close[knifeblock_76,cupboard_117]=True
    close[knifeblock_76,kitchen_counter_119]=True
    close[knifeblock_76,sink_120]=True
    close[knifeblock_76,faucet_121]=True
    close[knifeblock_76,stovefan_125]=True
    close[knifeblock_76,oven_127]=True
    close[knifeblock_76,tray_128]=True
    close[knifeblock_76,walllamp_140]=True
    close[knifeblock_76,walllamp_141]=True
    close[pot_78,floor_46]=True
    close[pot_78,ceiling_55]=True
    close[pot_78,wall_64]=True
    close[pot_78,wall_67]=True
    close[pot_78,wall_68]=True
    close[pot_78,knifeblock_76]=True
    close[pot_78,cupboard_117]=True
    close[pot_78,cupboard_118]=True
    close[pot_78,kitchen_counter_119]=True
    close[pot_78,sink_120]=True
    close[pot_78,kitchen_counter_122]=True
    close[pot_78,stovefan_125]=True
    close[pot_78,oven_127]=True
    close[pot_78,tray_128]=True
    close[pot_78,toaster_132]=True
    close[pot_78,walllamp_141]=True
    close[trashcan_99,vacuum_cleaner_2139]=True
    close[trashcan_99,floor_50]=True
    close[trashcan_99,floor_51]=True
    close[trashcan_99,wall_65]=True
    close[trashcan_99,wall_68]=True
    close[trashcan_99,kitchen_counter_122]=True
    close[trashcan_99,dishwasher_129]=True
    close[trashcan_99,coffe_maker_130]=True
    close[trashcan_99,wall_246]=True
    close[trashcan_99,floor_262]=True
    close[trashcan_99,bookshelf_275]=True
    close[trashcan_99,food_onion_2009]=True
    close[trashcan_99,glue_2045]=True
    close[trashcan_99,food_orange_2061]=True
    close[mat_102,floor_42]=True
    close[mat_102,floor_43]=True
    close[mat_102,floor_44]=True
    close[mat_102,floor_46]=True
    close[mat_102,floor_47]=True
    close[mat_102,floor_48]=True
    close[mat_102,floor_49]=True
    close[mat_102,floor_50]=True
    close[mat_102,pillow_103]=True
    close[mat_102,pillow_104]=True
    close[mat_102,pillow_105]=True
    close[mat_102,pillow_106]=True
    close[mat_102,bench_113]=True
    close[mat_102,table_114]=True
    close[mat_102,bench_115]=True
    close[mat_102,lighter_2004]=True
    close[mat_102,lighter_2039]=True
    close[pillow_103,floor_46]=True
    close[pillow_103,floor_47]=True
    close[pillow_103,floor_50]=True
    close[pillow_103,floor_51]=True
    close[pillow_103,wall_68]=True
    close[pillow_103,mat_102]=True
    close[pillow_103,pillow_104]=True
    close[pillow_103,pillow_105]=True
    close[pillow_103,pillow_106]=True
    close[pillow_103,bench_113]=True
    close[pillow_103,table_114]=True
    close[pillow_103,bench_115]=True
    close[pillow_104,floor_44]=True
    close[pillow_104,floor_45]=True
    close[pillow_104,floor_46]=True
    close[pillow_104,floor_47]=True
    close[pillow_104,wall_67]=True
    close[pillow_104,mat_102]=True
    close[pillow_104,pillow_103]=True
    close[pillow_104,pillow_105]=True
    close[pillow_104,pillow_106]=True
    close[pillow_104,bench_113]=True
    close[pillow_104,table_114]=True
    close[pillow_104,bench_115]=True
    close[pillow_105,floor_47]=True
    close[pillow_105,floor_48]=True
    close[pillow_105,floor_49]=True
    close[pillow_105,floor_50]=True
    close[pillow_105,wall_69]=True
    close[pillow_105,mat_102]=True
    close[pillow_105,pillow_103]=True
    close[pillow_105,pillow_104]=True
    close[pillow_105,pillow_106]=True
    close[pillow_105,bench_113]=True
    close[pillow_105,table_114]=True
    close[pillow_105,bench_115]=True
    close[pillow_106,floor_42]=True
    close[pillow_106,floor_43]=True
    close[pillow_106,floor_44]=True
    close[pillow_106,floor_47]=True
    close[pillow_106,floor_48]=True
    close[pillow_106,wall_70]=True
    close[pillow_106,mat_102]=True
    close[pillow_106,pillow_103]=True
    close[pillow_106,pillow_104]=True
    close[pillow_106,pillow_105]=True
    close[pillow_106,bench_113]=True
    close[pillow_106,table_114]=True
    close[pillow_106,bench_115]=True
    close[pillow_107,floor_48]=True
    close[pillow_107,floor_49]=True
    close[pillow_107,wall_63]=True
    close[pillow_107,wall_69]=True
    close[pillow_107,phone_71]=True
    close[pillow_107,pillow_108]=True
    close[pillow_107,drawing_111]=True
    close[pillow_107,tvstand_116]=True
    close[pillow_108,wall_2]=True
    close[pillow_108,floor_12]=True
    close[pillow_108,doorjamb_37]=True
    close[pillow_108,door_38]=True
    close[pillow_108,light_39]=True
    close[pillow_108,floor_42]=True
    close[pillow_108,floor_43]=True
    close[pillow_108,floor_48]=True
    close[pillow_108,wall_63]=True
    close[pillow_108,wall_70]=True
    close[pillow_108,pillow_107]=True
    close[pillow_108,drawing_111]=True
    close[pillow_108,tvstand_116]=True
    close[drawing_110,door_38]=True
    close[drawing_110,ceiling_52]=True
    close[drawing_110,ceiling_53]=True
    close[drawing_110,wall_66]=True
    close[drawing_110,wall_70]=True
    close[drawing_110,bookshelf_124]=True
    close[drawing_110,wall_176]=True
    close[drawing_110,wall_179]=True
    close[drawing_110,ceiling_182]=True
    close[drawing_110,ceiling_183]=True
    close[drawing_110,bookshelf_196]=True
    close[drawing_110,light_212]=True
    close[drawing_110,photoframe_219]=True
    close[drawing_111,wall_2]=True
    close[drawing_111,light_39]=True
    close[drawing_111,floor_48]=True
    close[drawing_111,ceiling_57]=True
    close[drawing_111,wall_63]=True
    close[drawing_111,wall_69]=True
    close[drawing_111,wall_70]=True
    close[drawing_111,phone_71]=True
    close[drawing_111,pillow_107]=True
    close[drawing_111,pillow_108]=True
    close[drawing_111,tvstand_116]=True
    close[bench_113,floor_44]=True
    close[bench_113,floor_45]=True
    close[bench_113,floor_46]=True
    close[bench_113,floor_47]=True
    close[bench_113,floor_50]=True
    close[bench_113,floor_51]=True
    close[bench_113,wall_67]=True
    close[bench_113,wall_68]=True
    close[bench_113,mat_102]=True
    close[bench_113,pillow_103]=True
    close[bench_113,pillow_104]=True
    close[bench_113,pillow_105]=True
    close[bench_113,pillow_106]=True
    close[bench_113,table_114]=True
    close[bench_113,bench_115]=True
    close[table_114,food_bread_2084]=True
    close[table_114,dry_pasta_2114]=True
    close[table_114,milk_2115]=True
    close[table_114,clothes_hat_2117]=True
    close[table_114,clothes_gloves_2118]=True
    close[table_114,knife_2122]=True
    close[table_114,cup_2132]=True
    close[table_114,cup_2133]=True
    close[table_114,cup_2134]=True
    close[table_114,floor_44]=True
    close[table_114,floor_47]=True
    close[table_114,floor_48]=True
    close[table_114,floor_50]=True
    close[table_114,mat_102]=True
    close[table_114,pillow_103]=True
    close[table_114,pillow_104]=True
    close[table_114,pillow_105]=True
    close[table_114,pillow_106]=True
    close[table_114,bench_113]=True
    close[table_114,bench_115]=True
    close[table_114,table_cloth_2005]=True
    close[table_114,food_food_2021]=True
    close[table_114,box_2038]=True
    close[table_114,cup_2049]=True
    close[table_114,check_2058]=True
    close[bench_115,floor_42]=True
    close[bench_115,floor_43]=True
    close[bench_115,floor_44]=True
    close[bench_115,floor_47]=True
    close[bench_115,floor_48]=True
    close[bench_115,floor_49]=True
    close[bench_115,floor_50]=True
    close[bench_115,wall_69]=True
    close[bench_115,wall_70]=True
    close[bench_115,mat_102]=True
    close[bench_115,pillow_103]=True
    close[bench_115,pillow_104]=True
    close[bench_115,pillow_105]=True
    close[bench_115,pillow_106]=True
    close[bench_115,bench_113]=True
    close[bench_115,table_114]=True
    close[tvstand_116,wall_2]=True
    close[tvstand_116,floor_12]=True
    close[tvstand_116,door_38]=True
    close[tvstand_116,light_39]=True
    close[tvstand_116,floor_42]=True
    close[tvstand_116,floor_43]=True
    close[tvstand_116,floor_48]=True
    close[tvstand_116,floor_49]=True
    close[tvstand_116,wall_63]=True
    close[tvstand_116,wall_69]=True
    close[tvstand_116,wall_70]=True
    close[tvstand_116,phone_71]=True
    close[tvstand_116,pillow_107]=True
    close[tvstand_116,pillow_108]=True
    close[tvstand_116,drawing_111]=True
    close[cupboard_117,ceiling_54]=True
    close[cupboard_117,ceiling_55]=True
    close[cupboard_117,wall_64]=True
    close[cupboard_117,wall_67]=True
    close[cupboard_117,knifeblock_76]=True
    close[cupboard_117,pot_78]=True
    close[cupboard_117,kitchen_counter_119]=True
    close[cupboard_117,sink_120]=True
    close[cupboard_117,faucet_121]=True
    close[cupboard_117,kitchen_counter_123]=True
    close[cupboard_117,stovefan_125]=True
    close[cupboard_117,oven_127]=True
    close[cupboard_117,tray_128]=True
    close[cupboard_117,walllamp_140]=True
    close[cupboard_117,walllamp_141]=True
    close[cupboard_117,coffee_filter_2053]=True
    close[cupboard_118,ceiling_55]=True
    close[cupboard_118,ceiling_60]=True
    close[cupboard_118,wall_64]=True
    close[cupboard_118,wall_68]=True
    close[cupboard_118,pot_78]=True
    close[cupboard_118,kitchen_counter_122]=True
    close[cupboard_118,stovefan_125]=True
    close[cupboard_118,oven_127]=True
    close[cupboard_118,tray_128]=True
    close[cupboard_118,dishwasher_129]=True
    close[cupboard_118,coffe_maker_130]=True
    close[cupboard_118,toaster_132]=True
    close[cupboard_118,microwave_135]=True
    close[cupboard_118,walllamp_139]=True
    close[cupboard_118,walllamp_141]=True
    close[cupboard_118,knife_2037]=True
    close[cupboard_118,tea_2066]=True
    close[cupboard_118,food_peanut_butter_2077]=True
    close[kitchen_counter_119,cutting_board_2123]=True
    close[kitchen_counter_119,stove_2135]=True
    close[kitchen_counter_119,pot_2138]=True
    close[kitchen_counter_119,bowl_2140]=True
    close[kitchen_counter_119,bowl_2141]=True
    close[kitchen_counter_119,bowl_2142]=True
    close[kitchen_counter_119,fork_2150]=True
    close[kitchen_counter_119,fork_2151]=True
    close[kitchen_counter_119,plate_2152]=True
    close[kitchen_counter_119,floor_45]=True
    close[kitchen_counter_119,floor_46]=True
    close[kitchen_counter_119,wall_64]=True
    close[kitchen_counter_119,wall_67]=True
    close[kitchen_counter_119,knifeblock_76]=True
    close[kitchen_counter_119,pot_78]=True
    close[kitchen_counter_119,cupboard_117]=True
    close[kitchen_counter_119,sink_120]=True
    close[kitchen_counter_119,faucet_121]=True
    close[kitchen_counter_119,kitchen_counter_123]=True
    close[kitchen_counter_119,stovefan_125]=True
    close[kitchen_counter_119,oven_127]=True
    close[kitchen_counter_119,tray_128]=True
    close[kitchen_counter_119,walllamp_140]=True
    close[kitchen_counter_119,walllamp_141]=True
    close[kitchen_counter_119,desk_193]=True
    close[kitchen_counter_119,cpuscreen_210]=True
    close[kitchen_counter_119,food_salt_2041]=True
    close[sink_120,basket_for_clothes_2078]=True
    close[sink_120,washing_machine_2079]=True
    close[sink_120,soap_2126]=True
    close[sink_120,floor_45]=True
    close[sink_120,floor_46]=True
    close[sink_120,wall_64]=True
    close[sink_120,wall_67]=True
    close[sink_120,knifeblock_76]=True
    close[sink_120,pot_78]=True
    close[sink_120,cupboard_117]=True
    close[sink_120,kitchen_counter_119]=True
    close[sink_120,faucet_121]=True
    close[sink_120,kitchen_counter_123]=True
    close[sink_120,walllamp_140]=True
    close[sink_120,soap_2010]=True
    close[sink_120,ice_2024]=True
    close[faucet_121,floor_45]=True
    close[faucet_121,floor_46]=True
    close[faucet_121,ceiling_54]=True
    close[faucet_121,wall_64]=True
    close[faucet_121,wall_67]=True
    close[faucet_121,knifeblock_76]=True
    close[faucet_121,cupboard_117]=True
    close[faucet_121,kitchen_counter_119]=True
    close[faucet_121,sink_120]=True
    close[faucet_121,oven_127]=True
    close[faucet_121,walllamp_140]=True
    close[kitchen_counter_122,spectacles_2153]=True
    close[kitchen_counter_122,fryingpan_2154]=True
    close[kitchen_counter_122,floor_46]=True
    close[kitchen_counter_122,floor_51]=True
    close[kitchen_counter_122,wall_64]=True
    close[kitchen_counter_122,wall_68]=True
    close[kitchen_counter_122,pot_78]=True
    close[kitchen_counter_122,trashcan_99]=True
    close[kitchen_counter_122,cupboard_118]=True
    close[kitchen_counter_122,stovefan_125]=True
    close[kitchen_counter_122,oven_127]=True
    close[kitchen_counter_122,tray_128]=True
    close[kitchen_counter_122,dishwasher_129]=True
    close[kitchen_counter_122,coffe_maker_130]=True
    close[kitchen_counter_122,toaster_132]=True
    close[kitchen_counter_122,microwave_135]=True
    close[kitchen_counter_122,walllamp_139]=True
    close[kitchen_counter_122,walllamp_141]=True
    close[kitchen_counter_123,oil_2149]=True
    close[kitchen_counter_123,floor_45]=True
    close[kitchen_counter_123,wall_67]=True
    close[kitchen_counter_123,cupboard_117]=True
    close[kitchen_counter_123,kitchen_counter_119]=True
    close[kitchen_counter_123,sink_120]=True
    close[kitchen_counter_123,floor_163]=True
    close[kitchen_counter_123,floor_164]=True
    close[kitchen_counter_123,wall_175]=True
    close[kitchen_counter_123,desk_193]=True
    close[kitchen_counter_123,cpuscreen_210]=True
    close[kitchen_counter_123,keyboard_211]=True
    close[kitchen_counter_123,food_orange_2027]=True
    close[kitchen_counter_123,knife_2035]=True
    close[kitchen_counter_123,food_kiwi_2054]=True
    close[kitchen_counter_123,tray_2068]=True
    close[bookshelf_124,book_2136]=True
    close[bookshelf_124,book_2137]=True
    close[bookshelf_124,doorjamb_37]=True
    close[bookshelf_124,door_38]=True
    close[bookshelf_124,floor_42]=True
    close[bookshelf_124,floor_43]=True
    close[bookshelf_124,floor_44]=True
    close[bookshelf_124,wall_66]=True
    close[bookshelf_124,wall_70]=True
    close[bookshelf_124,powersocket_72]=True
    close[bookshelf_124,drawing_110]=True
    close[bookshelf_124,floor_169]=True
    close[bookshelf_124,floor_170]=True
    close[bookshelf_124,wall_176]=True
    close[bookshelf_124,wall_179]=True
    close[bookshelf_124,bookshelf_196]=True
    close[bookshelf_124,light_212]=True
    close[bookshelf_124,photoframe_219]=True
    close[bookshelf_124,envelope_2055]=True
    close[stovefan_125,ceiling_54]=True
    close[stovefan_125,ceiling_55]=True
    close[stovefan_125,ceiling_60]=True
    close[stovefan_125,wall_64]=True
    close[stovefan_125,wall_67]=True
    close[stovefan_125,wall_68]=True
    close[stovefan_125,knifeblock_76]=True
    close[stovefan_125,pot_78]=True
    close[stovefan_125,cupboard_117]=True
    close[stovefan_125,cupboard_118]=True
    close[stovefan_125,kitchen_counter_119]=True
    close[stovefan_125,kitchen_counter_122]=True
    close[stovefan_125,oven_127]=True
    close[stovefan_125,tray_128]=True
    close[stovefan_125,toaster_132]=True
    close[stovefan_125,walllamp_141]=True
    close[fridge_126,basket_for_clothes_2078]=True
    close[fridge_126,washing_machine_2079]=True
    close[fridge_126,food_steak_2080]=True
    close[fridge_126,food_apple_2081]=True
    close[fridge_126,food_bacon_2082]=True
    close[fridge_126,food_banana_2083]=True
    close[fridge_126,food_cake_2085]=True
    close[fridge_126,food_carrot_2086]=True
    close[fridge_126,food_cereal_2087]=True
    close[fridge_126,food_cheese_2088]=True
    close[fridge_126,food_chicken_2089]=True
    close[fridge_126,food_dessert_2090]=True
    close[fridge_126,food_donut_2091]=True
    close[fridge_126,food_egg_2092]=True
    close[fridge_126,food_fish_2093]=True
    close[fridge_126,food_food_2094]=True
    close[fridge_126,food_fruit_2095]=True
    close[fridge_126,food_hamburger_2096]=True
    close[fridge_126,food_ice_cream_2097]=True
    close[fridge_126,food_jam_2098]=True
    close[fridge_126,food_kiwi_2099]=True
    close[fridge_126,food_lemon_2100]=True
    close[fridge_126,food_noodles_2101]=True
    close[fridge_126,food_oatmeal_2102]=True
    close[fridge_126,food_orange_2103]=True
    close[fridge_126,food_onion_2104]=True
    close[fridge_126,food_peanut_butter_2105]=True
    close[fridge_126,food_pizza_2106]=True
    close[fridge_126,food_potato_2107]=True
    close[fridge_126,food_rice_2108]=True
    close[fridge_126,food_salt_2109]=True
    close[fridge_126,food_snack_2110]=True
    close[fridge_126,food_sugar_2111]=True
    close[fridge_126,food_turkey_2112]=True
    close[fridge_126,food_vegetable_2113]=True
    close[fridge_126,sauce_2148]=True
    close[fridge_126,floor_44]=True
    close[fridge_126,floor_45]=True
    close[fridge_126,ceiling_53]=True
    close[fridge_126,ceiling_54]=True
    close[fridge_126,door_61]=True
    close[fridge_126,wall_66]=True
    close[fridge_126,wall_67]=True
    close[fridge_126,powersocket_72]=True
    close[fridge_126,light_73]=True
    close[fridge_126,ceilinglamp_137]=True
    close[fridge_126,floor_163]=True
    close[fridge_126,floor_164]=True
    close[fridge_126,floor_169]=True
    close[fridge_126,wall_175]=True
    close[fridge_126,wall_179]=True
    close[fridge_126,doorjamb_190]=True
    close[fridge_126,desk_193]=True
    close[fridge_126,computer_209]=True
    close[fridge_126,cpuscreen_210]=True
    close[fridge_126,keyboard_211]=True
    close[fridge_126,light_212]=True
    close[fridge_126,mouse_213]=True
    close[fridge_126,mousepad_214]=True
    close[fridge_126,food_food_1000]=True
    close[fridge_126,food_food_2001]=True
    close[fridge_126,food_food_2046]=True
    close[fridge_126,food_onion_2048]=True
    close[fridge_126,food_food_2073]=True
    close[oven_127,floor_46]=True
    close[oven_127,floor_51]=True
    close[oven_127,ceiling_55]=True
    close[oven_127,wall_64]=True
    close[oven_127,wall_67]=True
    close[oven_127,wall_68]=True
    close[oven_127,knifeblock_76]=True
    close[oven_127,pot_78]=True
    close[oven_127,cupboard_117]=True
    close[oven_127,cupboard_118]=True
    close[oven_127,kitchen_counter_119]=True
    close[oven_127,faucet_121]=True
    close[oven_127,kitchen_counter_122]=True
    close[oven_127,stovefan_125]=True
    close[oven_127,tray_128]=True
    close[oven_127,toaster_132]=True
    close[oven_127,walllamp_141]=True
    close[oven_127,oil_2013]=True
    close[oven_127,food_carrot_2015]=True
    close[oven_127,food_food_2064]=True
    close[oven_127,food_cheese_2072]=True
    close[tray_128,floor_46]=True
    close[tray_128,floor_51]=True
    close[tray_128,wall_64]=True
    close[tray_128,wall_67]=True
    close[tray_128,wall_68]=True
    close[tray_128,knifeblock_76]=True
    close[tray_128,pot_78]=True
    close[tray_128,cupboard_117]=True
    close[tray_128,cupboard_118]=True
    close[tray_128,kitchen_counter_119]=True
    close[tray_128,kitchen_counter_122]=True
    close[tray_128,stovefan_125]=True
    close[tray_128,oven_127]=True
    close[tray_128,toaster_132]=True
    close[tray_128,walllamp_141]=True
    close[dishwasher_129,floor_46]=True
    close[dishwasher_129,floor_51]=True
    close[dishwasher_129,wall_64]=True
    close[dishwasher_129,wall_68]=True
    close[dishwasher_129,trashcan_99]=True
    close[dishwasher_129,cupboard_118]=True
    close[dishwasher_129,kitchen_counter_122]=True
    close[dishwasher_129,coffe_maker_130]=True
    close[dishwasher_129,toaster_132]=True
    close[dishwasher_129,microwave_135]=True
    close[dishwasher_129,walllamp_139]=True
    close[dishwasher_129,detergent_2011]=True
    close[dishwasher_129,measuring_cup_2012]=True
    close[coffe_maker_130,floor_51]=True
    close[coffe_maker_130,ceiling_60]=True
    close[coffe_maker_130,wall_68]=True
    close[coffe_maker_130,trashcan_99]=True
    close[coffe_maker_130,cupboard_118]=True
    close[coffe_maker_130,kitchen_counter_122]=True
    close[coffe_maker_130,dishwasher_129]=True
    close[coffe_maker_130,toaster_132]=True
    close[coffe_maker_130,microwave_135]=True
    close[coffe_maker_130,walllamp_139]=True
    close[coffe_maker_130,coffee_filter_2065]=True
    close[toaster_132,floor_46]=True
    close[toaster_132,floor_51]=True
    close[toaster_132,ceiling_55]=True
    close[toaster_132,ceiling_60]=True
    close[toaster_132,wall_64]=True
    close[toaster_132,wall_68]=True
    close[toaster_132,pot_78]=True
    close[toaster_132,cupboard_118]=True
    close[toaster_132,kitchen_counter_122]=True
    close[toaster_132,stovefan_125]=True
    close[toaster_132,oven_127]=True
    close[toaster_132,tray_128]=True
    close[toaster_132,dishwasher_129]=True
    close[toaster_132,coffe_maker_130]=True
    close[toaster_132,microwave_135]=True
    close[toaster_132,walllamp_139]=True
    close[toaster_132,walllamp_141]=True
    close[microwave_135,floor_51]=True
    close[microwave_135,ceiling_60]=True
    close[microwave_135,wall_64]=True
    close[microwave_135,wall_68]=True
    close[microwave_135,cupboard_118]=True
    close[microwave_135,kitchen_counter_122]=True
    close[microwave_135,dishwasher_129]=True
    close[microwave_135,coffe_maker_130]=True
    close[microwave_135,toaster_132]=True
    close[microwave_135,walllamp_139]=True
    close[microwave_135,pot_2040]=True
    close[ceilinglamp_137,ceiling_52]=True
    close[ceilinglamp_137,ceiling_53]=True
    close[ceilinglamp_137,ceiling_54]=True
    close[ceilinglamp_137,ceiling_55]=True
    close[ceilinglamp_137,ceiling_56]=True
    close[ceilinglamp_137,ceiling_57]=True
    close[ceilinglamp_137,wall_67]=True
    close[ceilinglamp_137,wall_70]=True
    close[ceilinglamp_137,fridge_126]=True
    close[ceilinglamp_138,ceiling_55]=True
    close[ceilinglamp_138,ceiling_56]=True
    close[ceilinglamp_138,ceiling_57]=True
    close[ceilinglamp_138,ceiling_58]=True
    close[ceilinglamp_138,ceiling_59]=True
    close[ceilinglamp_138,ceiling_60]=True
    close[ceilinglamp_138,wall_68]=True
    close[ceilinglamp_138,wall_69]=True
    close[walllamp_139,ceiling_55]=True
    close[walllamp_139,ceiling_60]=True
    close[walllamp_139,wall_64]=True
    close[walllamp_139,wall_68]=True
    close[walllamp_139,cupboard_118]=True
    close[walllamp_139,kitchen_counter_122]=True
    close[walllamp_139,dishwasher_129]=True
    close[walllamp_139,coffe_maker_130]=True
    close[walllamp_139,toaster_132]=True
    close[walllamp_139,microwave_135]=True
    close[walllamp_140,ceiling_54]=True
    close[walllamp_140,ceiling_55]=True
    close[walllamp_140,wall_64]=True
    close[walllamp_140,wall_67]=True
    close[walllamp_140,knifeblock_76]=True
    close[walllamp_140,cupboard_117]=True
    close[walllamp_140,kitchen_counter_119]=True
    close[walllamp_140,sink_120]=True
    close[walllamp_140,faucet_121]=True
    close[walllamp_141,ceiling_55]=True
    close[walllamp_141,ceiling_60]=True
    close[walllamp_141,wall_64]=True
    close[walllamp_141,wall_67]=True
    close[walllamp_141,wall_68]=True
    close[walllamp_141,knifeblock_76]=True
    close[walllamp_141,pot_78]=True
    close[walllamp_141,cupboard_117]=True
    close[walllamp_141,cupboard_118]=True
    close[walllamp_141,kitchen_counter_119]=True
    close[walllamp_141,kitchen_counter_122]=True
    close[walllamp_141,stovefan_125]=True
    close[walllamp_141,oven_127]=True
    close[walllamp_141,tray_128]=True
    close[walllamp_141,toaster_132]=True
    close[floor_163,floor_45]=True
    close[floor_163,door_61]=True
    close[floor_163,wall_67]=True
    close[floor_163,light_73]=True
    close[floor_163,kitchen_counter_123]=True
    close[floor_163,fridge_126]=True
    close[floor_163,floor_164]=True
    close[floor_163,floor_165]=True
    close[floor_163,floor_169]=True
    close[floor_163,wall_175]=True
    close[floor_163,desk_193]=True
    close[floor_163,chair_194]=True
    close[floor_163,nightstand_195]=True
    close[floor_163,computer_209]=True
    close[floor_163,cpuscreen_210]=True
    close[floor_163,keyboard_211]=True
    close[floor_163,mouse_213]=True
    close[floor_163,mousepad_214]=True
    close[floor_164,floor_45]=True
    close[floor_164,door_61]=True
    close[floor_164,wall_67]=True
    close[floor_164,light_73]=True
    close[floor_164,kitchen_counter_123]=True
    close[floor_164,fridge_126]=True
    close[floor_164,floor_163]=True
    close[floor_164,floor_165]=True
    close[floor_164,floor_169]=True
    close[floor_164,wall_175]=True
    close[floor_164,desk_193]=True
    close[floor_164,chair_194]=True
    close[floor_164,nightstand_195]=True
    close[floor_164,computer_209]=True
    close[floor_164,cpuscreen_210]=True
    close[floor_164,keyboard_211]=True
    close[floor_164,mouse_213]=True
    close[floor_164,mousepad_214]=True
    close[floor_165,floor_163]=True
    close[floor_165,floor_164]=True
    close[floor_165,floor_166]=True
    close[floor_165,floor_168]=True
    close[floor_165,wall_173]=True
    close[floor_165,wall_175]=True
    close[floor_165,wall_178]=True
    close[floor_165,chair_194]=True
    close[floor_165,nightstand_195]=True
    close[floor_165,bed_197]=True
    close[floor_165,drawing_201]=True
    close[floor_165,pillow_207]=True
    close[floor_165,pillow_208]=True
    close[floor_165,tablelamp_239]=True
    close[floor_166,floor_165]=True
    close[floor_166,floor_167]=True
    close[floor_166,wall_178]=True
    close[floor_166,nightstand_192]=True
    close[floor_166,nightstand_195]=True
    close[floor_166,bed_197]=True
    close[floor_166,drawing_201]=True
    close[floor_166,pillow_207]=True
    close[floor_166,pillow_208]=True
    close[floor_166,tablelamp_238]=True
    close[floor_166,tablelamp_239]=True
    close[floor_167,floor_166]=True
    close[floor_167,floor_168]=True
    close[floor_167,floor_172]=True
    close[floor_167,wall_177]=True
    close[floor_167,wall_178]=True
    close[floor_167,wall_180]=True
    close[floor_167,window_191]=True
    close[floor_167,bed_197]=True
    close[floor_167,table_199]=True
    close[floor_167,mat_203]=True
    close[floor_167,curtain_204]=True
    close[floor_167,curtain_205]=True
    close[floor_167,curtain_206]=True
    close[floor_168,floor_165]=True
    close[floor_168,floor_167]=True
    close[floor_168,floor_169]=True
    close[floor_168,floor_171]=True
    close[floor_168,chair_194]=True
    close[floor_168,bed_197]=True
    close[floor_168,table_199]=True
    close[floor_168,mat_203]=True
    close[floor_169,floor_44]=True
    close[floor_169,door_61]=True
    close[floor_169,wall_66]=True
    close[floor_169,powersocket_72]=True
    close[floor_169,light_73]=True
    close[floor_169,bookshelf_124]=True
    close[floor_169,fridge_126]=True
    close[floor_169,floor_163]=True
    close[floor_169,floor_164]=True
    close[floor_169,floor_168]=True
    close[floor_169,floor_170]=True
    close[floor_169,wall_175]=True
    close[floor_169,wall_176]=True
    close[floor_169,wall_179]=True
    close[floor_169,doorjamb_190]=True
    close[floor_169,desk_193]=True
    close[floor_169,chair_194]=True
    close[floor_169,bookshelf_196]=True
    close[floor_169,mat_203]=True
    close[floor_169,computer_209]=True
    close[floor_169,keyboard_211]=True
    close[floor_169,light_212]=True
    close[floor_169,mouse_213]=True
    close[floor_169,mousepad_214]=True
    close[floor_170,wall_5]=True
    close[floor_170,floor_13]=True
    close[floor_170,toilet_15]=True
    close[floor_170,shower_16]=True
    close[floor_170,shower_21]=True
    close[floor_170,door_38]=True
    close[floor_170,floor_42]=True
    close[floor_170,floor_43]=True
    close[floor_170,door_61]=True
    close[floor_170,wall_70]=True
    close[floor_170,powersocket_72]=True
    close[floor_170,bookshelf_124]=True
    close[floor_170,floor_169]=True
    close[floor_170,floor_171]=True
    close[floor_170,wall_176]=True
    close[floor_170,bookshelf_196]=True
    close[floor_170,filing_cabinet_200]=True
    close[floor_170,mat_203]=True
    close[floor_170,light_212]=True
    close[floor_170,photoframe_219]=True
    close[floor_171,floor_168]=True
    close[floor_171,floor_170]=True
    close[floor_171,floor_172]=True
    close[floor_171,wall_174]=True
    close[floor_171,wall_176]=True
    close[floor_171,wall_177]=True
    close[floor_171,couch_198]=True
    close[floor_171,table_199]=True
    close[floor_171,filing_cabinet_200]=True
    close[floor_171,mat_203]=True
    close[floor_172,floor_167]=True
    close[floor_172,floor_171]=True
    close[floor_172,wall_177]=True
    close[floor_172,couch_198]=True
    close[floor_172,table_199]=True
    close[floor_172,mat_203]=True
    close[wall_173,floor_165]=True
    close[wall_173,wall_175]=True
    close[wall_173,wall_178]=True
    close[wall_173,ceiling_186]=True
    close[wall_173,nightstand_195]=True
    close[wall_173,bed_197]=True
    close[wall_173,drawing_201]=True
    close[wall_173,pillow_207]=True
    close[wall_173,pillow_208]=True
    close[wall_173,tablelamp_239]=True
    close[wall_174,wall_5]=True
    close[wall_174,shower_21]=True
    close[wall_174,floor_171]=True
    close[wall_174,wall_176]=True
    close[wall_174,wall_177]=True
    close[wall_174,ceiling_184]=True
    close[wall_174,couch_198]=True
    close[wall_174,filing_cabinet_200]=True
    close[wall_174,drawing_202]=True
    close[wall_174,mat_203]=True
    close[wall_175,floor_45]=True
    close[wall_175,ceiling_54]=True
    close[wall_175,door_61]=True
    close[wall_175,wall_66]=True
    close[wall_175,wall_67]=True
    close[wall_175,light_73]=True
    close[wall_175,kitchen_counter_123]=True
    close[wall_175,fridge_126]=True
    close[wall_175,floor_163]=True
    close[wall_175,floor_164]=True
    close[wall_175,floor_165]=True
    close[wall_175,floor_169]=True
    close[wall_175,wall_173]=True
    close[wall_175,wall_179]=True
    close[wall_175,ceiling_181]=True
    close[wall_175,ceiling_182]=True
    close[wall_175,ceiling_186]=True
    close[wall_175,doorjamb_190]=True
    close[wall_175,desk_193]=True
    close[wall_175,chair_194]=True
    close[wall_175,nightstand_195]=True
    close[wall_175,computer_209]=True
    close[wall_175,cpuscreen_210]=True
    close[wall_175,keyboard_211]=True
    close[wall_175,mouse_213]=True
    close[wall_175,mousepad_214]=True
    close[wall_175,tablelamp_239]=True
    close[wall_176,wall_5]=True
    close[wall_176,ceiling_8]=True
    close[wall_176,floor_13]=True
    close[wall_176,toilet_15]=True
    close[wall_176,shower_16]=True
    close[wall_176,shower_21]=True
    close[wall_176,doorjamb_37]=True
    close[wall_176,door_38]=True
    close[wall_176,floor_42]=True
    close[wall_176,floor_43]=True
    close[wall_176,ceiling_52]=True
    close[wall_176,door_61]=True
    close[wall_176,wall_66]=True
    close[wall_176,wall_70]=True
    close[wall_176,powersocket_72]=True
    close[wall_176,drawing_110]=True
    close[wall_176,bookshelf_124]=True
    close[wall_176,floor_169]=True
    close[wall_176,floor_170]=True
    close[wall_176,floor_171]=True
    close[wall_176,wall_174]=True
    close[wall_176,wall_179]=True
    close[wall_176,ceiling_182]=True
    close[wall_176,ceiling_183]=True
    close[wall_176,ceiling_184]=True
    close[wall_176,doorjamb_190]=True
    close[wall_176,bookshelf_196]=True
    close[wall_176,filing_cabinet_200]=True
    close[wall_176,drawing_202]=True
    close[wall_176,light_212]=True
    close[wall_176,photoframe_219]=True
    close[wall_176,ceilinglamp_237]=True
    close[wall_177,floor_167]=True
    close[wall_177,floor_171]=True
    close[wall_177,floor_172]=True
    close[wall_177,wall_174]=True
    close[wall_177,wall_180]=True
    close[wall_177,ceiling_184]=True
    close[wall_177,ceiling_188]=True
    close[wall_177,ceiling_189]=True
    close[wall_177,window_191]=True
    close[wall_177,couch_198]=True
    close[wall_177,table_199]=True
    close[wall_177,mat_203]=True
    close[wall_177,curtain_206]=True
    close[wall_178,floor_165]=True
    close[wall_178,floor_166]=True
    close[wall_178,floor_167]=True
    close[wall_178,wall_173]=True
    close[wall_178,wall_180]=True
    close[wall_178,ceiling_186]=True
    close[wall_178,ceiling_187]=True
    close[wall_178,ceiling_188]=True
    close[wall_178,window_191]=True
    close[wall_178,nightstand_192]=True
    close[wall_178,nightstand_195]=True
    close[wall_178,bed_197]=True
    close[wall_178,drawing_201]=True
    close[wall_178,curtain_204]=True
    close[wall_178,curtain_205]=True
    close[wall_178,pillow_207]=True
    close[wall_178,pillow_208]=True
    close[wall_178,tablelamp_238]=True
    close[wall_178,tablelamp_239]=True
    close[wall_179,floor_44]=True
    close[wall_179,ceiling_53]=True
    close[wall_179,door_61]=True
    close[wall_179,wall_66]=True
    close[wall_179,wall_67]=True
    close[wall_179,wall_70]=True
    close[wall_179,powersocket_72]=True
    close[wall_179,light_73]=True
    close[wall_179,drawing_110]=True
    close[wall_179,bookshelf_124]=True
    close[wall_179,fridge_126]=True
    close[wall_179,floor_169]=True
    close[wall_179,wall_175]=True
    close[wall_179,wall_176]=True
    close[wall_179,ceiling_182]=True
    close[wall_179,doorjamb_190]=True
    close[wall_179,desk_193]=True
    close[wall_179,bookshelf_196]=True
    close[wall_179,computer_209]=True
    close[wall_179,cpuscreen_210]=True
    close[wall_179,keyboard_211]=True
    close[wall_179,light_212]=True
    close[wall_179,mouse_213]=True
    close[wall_179,mousepad_214]=True
    close[wall_180,floor_167]=True
    close[wall_180,wall_177]=True
    close[wall_180,wall_178]=True
    close[wall_180,ceiling_188]=True
    close[wall_180,window_191]=True
    close[wall_180,mat_203]=True
    close[wall_180,curtain_204]=True
    close[wall_180,curtain_205]=True
    close[wall_180,curtain_206]=True
    close[ceiling_181,ceiling_54]=True
    close[ceiling_181,wall_67]=True
    close[ceiling_181,wall_175]=True
    close[ceiling_181,ceiling_182]=True
    close[ceiling_181,ceiling_186]=True
    close[ceiling_181,chair_194]=True
    close[ceiling_181,cpuscreen_210]=True
    close[ceiling_182,ceiling_53]=True
    close[ceiling_182,wall_66]=True
    close[ceiling_182,light_73]=True
    close[ceiling_182,drawing_110]=True
    close[ceiling_182,wall_175]=True
    close[ceiling_182,wall_176]=True
    close[ceiling_182,wall_179]=True
    close[ceiling_182,ceiling_181]=True
    close[ceiling_182,ceiling_183]=True
    close[ceiling_182,ceiling_185]=True
    close[ceiling_182,doorjamb_190]=True
    close[ceiling_182,bookshelf_196]=True
    close[ceiling_182,light_212]=True
    close[ceiling_182,ceilinglamp_237]=True
    close[ceiling_183,wall_5]=True
    close[ceiling_183,ceiling_8]=True
    close[ceiling_183,shower_16]=True
    close[ceiling_183,shower_21]=True
    close[ceiling_183,ceiling_52]=True
    close[ceiling_183,wall_70]=True
    close[ceiling_183,drawing_110]=True
    close[ceiling_183,wall_176]=True
    close[ceiling_183,ceiling_182]=True
    close[ceiling_183,ceiling_184]=True
    close[ceiling_183,bookshelf_196]=True
    close[ceiling_183,drawing_202]=True
    close[ceiling_183,light_212]=True
    close[ceiling_183,ceilinglamp_237]=True
    close[ceiling_184,wall_174]=True
    close[ceiling_184,wall_176]=True
    close[ceiling_184,wall_177]=True
    close[ceiling_184,ceiling_183]=True
    close[ceiling_184,ceiling_185]=True
    close[ceiling_184,ceiling_189]=True
    close[ceiling_184,drawing_202]=True
    close[ceiling_184,ceilinglamp_237]=True
    close[ceiling_185,ceiling_182]=True
    close[ceiling_185,ceiling_184]=True
    close[ceiling_185,ceiling_186]=True
    close[ceiling_185,ceiling_188]=True
    close[ceiling_185,ceilinglamp_237]=True
    close[ceiling_186,wall_173]=True
    close[ceiling_186,wall_175]=True
    close[ceiling_186,wall_178]=True
    close[ceiling_186,ceiling_181]=True
    close[ceiling_186,ceiling_185]=True
    close[ceiling_186,ceiling_187]=True
    close[ceiling_186,chair_194]=True
    close[ceiling_186,drawing_201]=True
    close[ceiling_187,wall_178]=True
    close[ceiling_187,ceiling_186]=True
    close[ceiling_187,ceiling_188]=True
    close[ceiling_187,drawing_201]=True
    close[ceiling_187,curtain_204]=True
    close[ceiling_187,curtain_205]=True
    close[ceiling_188,wall_177]=True
    close[ceiling_188,wall_178]=True
    close[ceiling_188,wall_180]=True
    close[ceiling_188,ceiling_185]=True
    close[ceiling_188,ceiling_187]=True
    close[ceiling_188,ceiling_189]=True
    close[ceiling_188,window_191]=True
    close[ceiling_188,curtain_204]=True
    close[ceiling_188,curtain_205]=True
    close[ceiling_188,curtain_206]=True
    close[ceiling_189,wall_177]=True
    close[ceiling_189,ceiling_184]=True
    close[ceiling_189,ceiling_188]=True
    close[ceiling_189,curtain_206]=True
    close[doorjamb_190,floor_44]=True
    close[doorjamb_190,ceiling_53]=True
    close[doorjamb_190,door_61]=True
    close[doorjamb_190,wall_66]=True
    close[doorjamb_190,wall_67]=True
    close[doorjamb_190,wall_70]=True
    close[doorjamb_190,powersocket_72]=True
    close[doorjamb_190,light_73]=True
    close[doorjamb_190,fridge_126]=True
    close[doorjamb_190,floor_169]=True
    close[doorjamb_190,wall_175]=True
    close[doorjamb_190,wall_176]=True
    close[doorjamb_190,wall_179]=True
    close[doorjamb_190,ceiling_182]=True
    close[doorjamb_190,desk_193]=True
    close[doorjamb_190,bookshelf_196]=True
    close[doorjamb_190,computer_209]=True
    close[doorjamb_190,light_212]=True
    close[doorjamb_190,mouse_213]=True
    close[doorjamb_190,mousepad_214]=True
    close[window_191,floor_167]=True
    close[window_191,wall_177]=True
    close[window_191,wall_178]=True
    close[window_191,wall_180]=True
    close[window_191,ceiling_188]=True
    close[window_191,mat_203]=True
    close[window_191,curtain_204]=True
    close[window_191,curtain_205]=True
    close[window_191,curtain_206]=True
    close[nightstand_192,floor_166]=True
    close[nightstand_192,wall_178]=True
    close[nightstand_192,bed_197]=True
    close[nightstand_192,drawing_201]=True
    close[nightstand_192,pillow_208]=True
    close[nightstand_192,tablelamp_238]=True
    close[desk_193,floor_44]=True
    close[desk_193,floor_45]=True
    close[desk_193,door_61]=True
    close[desk_193,wall_66]=True
    close[desk_193,wall_67]=True
    close[desk_193,light_73]=True
    close[desk_193,kitchen_counter_119]=True
    close[desk_193,kitchen_counter_123]=True
    close[desk_193,fridge_126]=True
    close[desk_193,floor_163]=True
    close[desk_193,floor_164]=True
    close[desk_193,floor_169]=True
    close[desk_193,wall_175]=True
    close[desk_193,wall_179]=True
    close[desk_193,doorjamb_190]=True
    close[desk_193,chair_194]=True
    close[desk_193,computer_209]=True
    close[desk_193,cpuscreen_210]=True
    close[desk_193,keyboard_211]=True
    close[desk_193,mouse_213]=True
    close[desk_193,mousepad_214]=True
    close[desk_193,check_2026]=True
    close[desk_193,laser_pointer_2034]=True
    close[chair_194,floor_163]=True
    close[chair_194,floor_164]=True
    close[chair_194,floor_165]=True
    close[chair_194,floor_168]=True
    close[chair_194,floor_169]=True
    close[chair_194,wall_175]=True
    close[chair_194,ceiling_181]=True
    close[chair_194,ceiling_186]=True
    close[chair_194,desk_193]=True
    close[chair_194,nightstand_195]=True
    close[chair_194,computer_209]=True
    close[chair_194,keyboard_211]=True
    close[chair_194,mouse_213]=True
    close[chair_194,mousepad_214]=True
    close[chair_194,tablelamp_239]=True
    close[nightstand_195,floor_163]=True
    close[nightstand_195,floor_164]=True
    close[nightstand_195,floor_165]=True
    close[nightstand_195,floor_166]=True
    close[nightstand_195,wall_173]=True
    close[nightstand_195,wall_175]=True
    close[nightstand_195,wall_178]=True
    close[nightstand_195,chair_194]=True
    close[nightstand_195,bed_197]=True
    close[nightstand_195,drawing_201]=True
    close[nightstand_195,pillow_207]=True
    close[nightstand_195,pillow_208]=True
    close[nightstand_195,tablelamp_239]=True
    close[bookshelf_196,toilet_15]=True
    close[bookshelf_196,shower_16]=True
    close[bookshelf_196,doorjamb_37]=True
    close[bookshelf_196,door_38]=True
    close[bookshelf_196,floor_42]=True
    close[bookshelf_196,floor_43]=True
    close[bookshelf_196,floor_44]=True
    close[bookshelf_196,ceiling_52]=True
    close[bookshelf_196,door_61]=True
    close[bookshelf_196,wall_66]=True
    close[bookshelf_196,wall_70]=True
    close[bookshelf_196,powersocket_72]=True
    close[bookshelf_196,drawing_110]=True
    close[bookshelf_196,bookshelf_124]=True
    close[bookshelf_196,floor_169]=True
    close[bookshelf_196,floor_170]=True
    close[bookshelf_196,wall_176]=True
    close[bookshelf_196,wall_179]=True
    close[bookshelf_196,ceiling_182]=True
    close[bookshelf_196,ceiling_183]=True
    close[bookshelf_196,doorjamb_190]=True
    close[bookshelf_196,filing_cabinet_200]=True
    close[bookshelf_196,light_212]=True
    close[bookshelf_196,photoframe_219]=True
    close[bookshelf_196,novel_2060]=True
    close[bed_197,clothes_dress_2116]=True
    close[bed_197,clothes_scarf_2120]=True
    close[bed_197,clothes_underwear_2121]=True
    close[bed_197,floor_165]=True
    close[bed_197,floor_166]=True
    close[bed_197,floor_167]=True
    close[bed_197,floor_168]=True
    close[bed_197,wall_173]=True
    close[bed_197,wall_178]=True
    close[bed_197,nightstand_192]=True
    close[bed_197,nightstand_195]=True
    close[bed_197,drawing_201]=True
    close[bed_197,pillow_207]=True
    close[bed_197,pillow_208]=True
    close[bed_197,tablelamp_238]=True
    close[bed_197,tablelamp_239]=True
    close[couch_198,clothes_jacket_2119]=True
    close[couch_198,floor_171]=True
    close[couch_198,floor_172]=True
    close[couch_198,wall_174]=True
    close[couch_198,wall_177]=True
    close[couch_198,table_199]=True
    close[couch_198,mat_203]=True
    close[couch_198,chair_2003]=True
    close[couch_198,phone_2016]=True
    close[couch_198,rag_2052]=True
    close[table_199,floor_167]=True
    close[table_199,floor_168]=True
    close[table_199,floor_171]=True
    close[table_199,floor_172]=True
    close[table_199,wall_177]=True
    close[table_199,couch_198]=True
    close[table_199,mat_203]=True
    close[table_199,wooden_spoon_2000]=True
    close[table_199,tea_bag_2023]=True
    close[filing_cabinet_200,wall_5]=True
    close[filing_cabinet_200,floor_13]=True
    close[filing_cabinet_200,toilet_15]=True
    close[filing_cabinet_200,shower_16]=True
    close[filing_cabinet_200,shower_21]=True
    close[filing_cabinet_200,wall_70]=True
    close[filing_cabinet_200,floor_170]=True
    close[filing_cabinet_200,floor_171]=True
    close[filing_cabinet_200,wall_174]=True
    close[filing_cabinet_200,wall_176]=True
    close[filing_cabinet_200,bookshelf_196]=True
    close[filing_cabinet_200,drawing_202]=True
    close[filing_cabinet_200,mat_203]=True
    close[filing_cabinet_200,photoframe_219]=True
    close[filing_cabinet_200,diary_2008]=True
    close[filing_cabinet_200,envelope_2018]=True
    close[filing_cabinet_200,rag_2025]=True
    close[filing_cabinet_200,cd_2030]=True
    close[filing_cabinet_200,scrabble_2031]=True
    close[filing_cabinet_200,after_shave_2042]=True
    close[filing_cabinet_200,homework_2047]=True
    close[filing_cabinet_200,stereo_2050]=True
    close[filing_cabinet_200,after_shave_2051]=True
    close[filing_cabinet_200,food_food_2074]=True
    close[drawing_201,floor_165]=True
    close[drawing_201,floor_166]=True
    close[drawing_201,wall_173]=True
    close[drawing_201,wall_178]=True
    close[drawing_201,ceiling_186]=True
    close[drawing_201,ceiling_187]=True
    close[drawing_201,nightstand_192]=True
    close[drawing_201,nightstand_195]=True
    close[drawing_201,bed_197]=True
    close[drawing_201,pillow_207]=True
    close[drawing_201,pillow_208]=True
    close[drawing_201,tablelamp_238]=True
    close[drawing_201,tablelamp_239]=True
    close[drawing_202,wall_5]=True
    close[drawing_202,ceiling_8]=True
    close[drawing_202,shower_21]=True
    close[drawing_202,wall_174]=True
    close[drawing_202,wall_176]=True
    close[drawing_202,ceiling_183]=True
    close[drawing_202,ceiling_184]=True
    close[drawing_202,filing_cabinet_200]=True
    close[mat_203,floor_167]=True
    close[mat_203,floor_168]=True
    close[mat_203,floor_169]=True
    close[mat_203,floor_170]=True
    close[mat_203,floor_171]=True
    close[mat_203,floor_172]=True
    close[mat_203,wall_174]=True
    close[mat_203,wall_177]=True
    close[mat_203,wall_180]=True
    close[mat_203,window_191]=True
    close[mat_203,couch_198]=True
    close[mat_203,table_199]=True
    close[mat_203,filing_cabinet_200]=True
    close[mat_203,curtain_204]=True
    close[mat_203,curtain_205]=True
    close[mat_203,curtain_206]=True
    close[mat_203,shoe_rack_2044]=True
    close[curtain_204,floor_167]=True
    close[curtain_204,wall_178]=True
    close[curtain_204,wall_180]=True
    close[curtain_204,ceiling_187]=True
    close[curtain_204,ceiling_188]=True
    close[curtain_204,window_191]=True
    close[curtain_204,mat_203]=True
    close[curtain_204,curtain_205]=True
    close[curtain_204,curtain_206]=True
    close[curtain_205,floor_167]=True
    close[curtain_205,wall_178]=True
    close[curtain_205,wall_180]=True
    close[curtain_205,ceiling_187]=True
    close[curtain_205,ceiling_188]=True
    close[curtain_205,window_191]=True
    close[curtain_205,mat_203]=True
    close[curtain_205,curtain_204]=True
    close[curtain_205,curtain_206]=True
    close[curtain_206,floor_167]=True
    close[curtain_206,wall_177]=True
    close[curtain_206,wall_180]=True
    close[curtain_206,ceiling_188]=True
    close[curtain_206,ceiling_189]=True
    close[curtain_206,window_191]=True
    close[curtain_206,mat_203]=True
    close[curtain_206,curtain_204]=True
    close[curtain_206,curtain_205]=True
    close[pillow_207,floor_165]=True
    close[pillow_207,floor_166]=True
    close[pillow_207,wall_173]=True
    close[pillow_207,wall_178]=True
    close[pillow_207,nightstand_195]=True
    close[pillow_207,bed_197]=True
    close[pillow_207,drawing_201]=True
    close[pillow_207,pillow_208]=True
    close[pillow_207,tablelamp_239]=True
    close[pillow_208,floor_165]=True
    close[pillow_208,floor_166]=True
    close[pillow_208,wall_173]=True
    close[pillow_208,wall_178]=True
    close[pillow_208,nightstand_192]=True
    close[pillow_208,nightstand_195]=True
    close[pillow_208,bed_197]=True
    close[pillow_208,drawing_201]=True
    close[pillow_208,pillow_207]=True
    close[pillow_208,tablelamp_238]=True
    close[pillow_208,tablelamp_239]=True
    close[computer_209,floor_44]=True
    close[computer_209,floor_45]=True
    close[computer_209,door_61]=True
    close[computer_209,wall_66]=True
    close[computer_209,wall_67]=True
    close[computer_209,light_73]=True
    close[computer_209,fridge_126]=True
    close[computer_209,floor_163]=True
    close[computer_209,floor_164]=True
    close[computer_209,floor_169]=True
    close[computer_209,wall_175]=True
    close[computer_209,wall_179]=True
    close[computer_209,doorjamb_190]=True
    close[computer_209,desk_193]=True
    close[computer_209,chair_194]=True
    close[computer_209,cpuscreen_210]=True
    close[computer_209,keyboard_211]=True
    close[computer_209,mouse_213]=True
    close[computer_209,mousepad_214]=True
    close[cpuscreen_210,floor_45]=True
    close[cpuscreen_210,ceiling_54]=True
    close[cpuscreen_210,wall_66]=True
    close[cpuscreen_210,wall_67]=True
    close[cpuscreen_210,light_73]=True
    close[cpuscreen_210,kitchen_counter_119]=True
    close[cpuscreen_210,kitchen_counter_123]=True
    close[cpuscreen_210,fridge_126]=True
    close[cpuscreen_210,floor_163]=True
    close[cpuscreen_210,floor_164]=True
    close[cpuscreen_210,wall_175]=True
    close[cpuscreen_210,wall_179]=True
    close[cpuscreen_210,ceiling_181]=True
    close[cpuscreen_210,desk_193]=True
    close[cpuscreen_210,computer_209]=True
    close[cpuscreen_210,keyboard_211]=True
    close[cpuscreen_210,mouse_213]=True
    close[cpuscreen_210,mousepad_214]=True
    close[keyboard_211,floor_45]=True
    close[keyboard_211,wall_66]=True
    close[keyboard_211,wall_67]=True
    close[keyboard_211,light_73]=True
    close[keyboard_211,kitchen_counter_123]=True
    close[keyboard_211,fridge_126]=True
    close[keyboard_211,floor_163]=True
    close[keyboard_211,floor_164]=True
    close[keyboard_211,floor_169]=True
    close[keyboard_211,wall_175]=True
    close[keyboard_211,wall_179]=True
    close[keyboard_211,desk_193]=True
    close[keyboard_211,chair_194]=True
    close[keyboard_211,computer_209]=True
    close[keyboard_211,cpuscreen_210]=True
    close[keyboard_211,mouse_213]=True
    close[keyboard_211,mousepad_214]=True
    close[light_212,floor_42]=True
    close[light_212,floor_43]=True
    close[light_212,floor_44]=True
    close[light_212,ceiling_52]=True
    close[light_212,ceiling_53]=True
    close[light_212,door_61]=True
    close[light_212,wall_66]=True
    close[light_212,wall_70]=True
    close[light_212,powersocket_72]=True
    close[light_212,light_73]=True
    close[light_212,drawing_110]=True
    close[light_212,bookshelf_124]=True
    close[light_212,fridge_126]=True
    close[light_212,floor_169]=True
    close[light_212,floor_170]=True
    close[light_212,wall_176]=True
    close[light_212,wall_179]=True
    close[light_212,ceiling_182]=True
    close[light_212,ceiling_183]=True
    close[light_212,doorjamb_190]=True
    close[light_212,bookshelf_196]=True
    close[mouse_213,floor_44]=True
    close[mouse_213,floor_45]=True
    close[mouse_213,door_61]=True
    close[mouse_213,wall_66]=True
    close[mouse_213,wall_67]=True
    close[mouse_213,light_73]=True
    close[mouse_213,fridge_126]=True
    close[mouse_213,floor_163]=True
    close[mouse_213,floor_164]=True
    close[mouse_213,floor_169]=True
    close[mouse_213,wall_175]=True
    close[mouse_213,wall_179]=True
    close[mouse_213,doorjamb_190]=True
    close[mouse_213,desk_193]=True
    close[mouse_213,chair_194]=True
    close[mouse_213,computer_209]=True
    close[mouse_213,cpuscreen_210]=True
    close[mouse_213,keyboard_211]=True
    close[mouse_213,mousepad_214]=True
    close[mousepad_214,floor_44]=True
    close[mousepad_214,floor_45]=True
    close[mousepad_214,door_61]=True
    close[mousepad_214,wall_66]=True
    close[mousepad_214,wall_67]=True
    close[mousepad_214,light_73]=True
    close[mousepad_214,fridge_126]=True
    close[mousepad_214,floor_163]=True
    close[mousepad_214,floor_164]=True
    close[mousepad_214,floor_169]=True
    close[mousepad_214,wall_175]=True
    close[mousepad_214,wall_179]=True
    close[mousepad_214,doorjamb_190]=True
    close[mousepad_214,desk_193]=True
    close[mousepad_214,chair_194]=True
    close[mousepad_214,computer_209]=True
    close[mousepad_214,cpuscreen_210]=True
    close[mousepad_214,keyboard_211]=True
    close[mousepad_214,mouse_213]=True
    close[photoframe_219,wall_2]=True
    close[photoframe_219,wall_5]=True
    close[photoframe_219,floor_12]=True
    close[photoframe_219,floor_13]=True
    close[photoframe_219,toilet_15]=True
    close[photoframe_219,shower_16]=True
    close[photoframe_219,shower_21]=True
    close[photoframe_219,doorjamb_37]=True
    close[photoframe_219,door_38]=True
    close[photoframe_219,floor_42]=True
    close[photoframe_219,floor_43]=True
    close[photoframe_219,wall_70]=True
    close[photoframe_219,drawing_110]=True
    close[photoframe_219,bookshelf_124]=True
    close[photoframe_219,floor_170]=True
    close[photoframe_219,wall_176]=True
    close[photoframe_219,bookshelf_196]=True
    close[photoframe_219,filing_cabinet_200]=True
    close[ceilinglamp_237,wall_176]=True
    close[ceilinglamp_237,ceiling_182]=True
    close[ceilinglamp_237,ceiling_183]=True
    close[ceilinglamp_237,ceiling_184]=True
    close[ceilinglamp_237,ceiling_185]=True
    close[tablelamp_238,floor_166]=True
    close[tablelamp_238,wall_178]=True
    close[tablelamp_238,nightstand_192]=True
    close[tablelamp_238,bed_197]=True
    close[tablelamp_238,drawing_201]=True
    close[tablelamp_238,pillow_208]=True
    close[tablelamp_239,floor_165]=True
    close[tablelamp_239,floor_166]=True
    close[tablelamp_239,wall_173]=True
    close[tablelamp_239,wall_175]=True
    close[tablelamp_239,wall_178]=True
    close[tablelamp_239,chair_194]=True
    close[tablelamp_239,nightstand_195]=True
    close[tablelamp_239,bed_197]=True
    close[tablelamp_239,drawing_201]=True
    close[tablelamp_239,pillow_207]=True
    close[tablelamp_239,pillow_208]=True
    close[wall_242,wall_247]=True
    close[wall_242,wall_248]=True
    close[wall_242,ceiling_255]=True
    close[wall_242,floor_265]=True
    close[wall_242,couch_269]=True
    close[wall_242,drawing_288]=True
    close[wall_242,walllamp_306]=True
    close[wall_242,walllamp_307]=True
    close[wall_243,wall_246]=True
    close[wall_243,wall_249]=True
    close[wall_243,ceiling_253]=True
    close[wall_243,floor_263]=True
    close[wall_243,desk_272]=True
    close[wall_243,computer_276]=True
    close[wall_243,cpuscreen_277]=True
    close[wall_243,keyboard_278]=True
    close[wall_243,mousepad_279]=True
    close[wall_243,mouse_280]=True
    close[wall_243,walllamp_304]=True
    close[wall_243,walllamp_305]=True
    close[wall_243,doorjamb_308]=True
    close[wall_244,floor_49]=True
    close[wall_244,ceiling_58]=True
    close[wall_244,door_62]=True
    close[wall_244,wall_65]=True
    close[wall_244,wall_69]=True
    close[wall_244,wall_246]=True
    close[wall_244,wall_247]=True
    close[wall_244,ceiling_251]=True
    close[wall_244,floor_261]=True
    close[wall_244,tvstand_273]=True
    close[wall_244,television_281]=True
    close[wall_244,powersocket_282]=True
    close[wall_244,light_283]=True
    close[wall_244,mat_284]=True
    close[wall_244,doorjamb_309]=True
    close[wall_245,wall_248]=True
    close[wall_245,wall_249]=True
    close[wall_245,ceiling_257]=True
    close[wall_245,floor_267]=True
    close[wall_245,couch_269]=True
    close[wall_245,dresser_274]=True
    close[wall_245,pillow_286]=True
    close[wall_245,pillow_287]=True
    close[wall_245,curtain_289]=True
    close[wall_245,curtain_290]=True
    close[wall_245,curtain_291]=True
    close[wall_245,hanger_292]=True
    close[wall_245,hanger_293]=True
    close[wall_245,hanger_294]=True
    close[wall_245,window_310]=True
    close[wall_246,floor_50]=True
    close[wall_246,ceiling_59]=True
    close[wall_246,door_62]=True
    close[wall_246,wall_65]=True
    close[wall_246,trashcan_99]=True
    close[wall_246,wall_243]=True
    close[wall_246,wall_244]=True
    close[wall_246,ceiling_251]=True
    close[wall_246,ceiling_252]=True
    close[wall_246,ceiling_253]=True
    close[wall_246,floor_261]=True
    close[wall_246,floor_262]=True
    close[wall_246,floor_263]=True
    close[wall_246,chair_271]=True
    close[wall_246,desk_272]=True
    close[wall_246,bookshelf_275]=True
    close[wall_246,computer_276]=True
    close[wall_246,cpuscreen_277]=True
    close[wall_246,keyboard_278]=True
    close[wall_246,mousepad_279]=True
    close[wall_246,mouse_280]=True
    close[wall_246,light_283]=True
    close[wall_246,mat_284]=True
    close[wall_246,walllamp_304]=True
    close[wall_246,doorjamb_309]=True
    close[wall_247,door_62]=True
    close[wall_247,wall_242]=True
    close[wall_247,wall_244]=True
    close[wall_247,ceiling_250]=True
    close[wall_247,ceiling_251]=True
    close[wall_247,ceiling_255]=True
    close[wall_247,floor_259]=True
    close[wall_247,floor_260]=True
    close[wall_247,floor_261]=True
    close[wall_247,floor_265]=True
    close[wall_247,tvstand_273]=True
    close[wall_247,television_281]=True
    close[wall_247,powersocket_282]=True
    close[wall_247,mat_284]=True
    close[wall_247,drawing_288]=True
    close[wall_247,walllamp_306]=True
    close[wall_247,doorjamb_309]=True
    close[wall_248,wall_242]=True
    close[wall_248,wall_245]=True
    close[wall_248,ceiling_255]=True
    close[wall_248,ceiling_256]=True
    close[wall_248,ceiling_257]=True
    close[wall_248,floor_265]=True
    close[wall_248,floor_266]=True
    close[wall_248,floor_267]=True
    close[wall_248,couch_269]=True
    close[wall_248,table_270]=True
    close[wall_248,orchid_285]=True
    close[wall_248,pillow_286]=True
    close[wall_248,pillow_287]=True
    close[wall_248,curtain_291]=True
    close[wall_248,walllamp_307]=True
    close[wall_248,window_310]=True
    close[wall_249,wall_243]=True
    close[wall_249,wall_245]=True
    close[wall_249,ceiling_253]=True
    close[wall_249,ceiling_257]=True
    close[wall_249,ceiling_258]=True
    close[wall_249,floor_263]=True
    close[wall_249,floor_267]=True
    close[wall_249,floor_268]=True
    close[wall_249,dresser_274]=True
    close[wall_249,computer_276]=True
    close[wall_249,mousepad_279]=True
    close[wall_249,mouse_280]=True
    close[wall_249,curtain_289]=True
    close[wall_249,curtain_290]=True
    close[wall_249,hanger_292]=True
    close[wall_249,hanger_293]=True
    close[wall_249,hanger_294]=True
    close[wall_249,walllamp_305]=True
    close[wall_249,doorjamb_308]=True
    close[wall_249,window_310]=True
    close[ceiling_250,wall_247]=True
    close[ceiling_250,ceiling_251]=True
    close[ceiling_250,ceiling_255]=True
    close[ceiling_250,television_281]=True
    close[ceiling_250,drawing_288]=True
    close[ceiling_250,walllamp_306]=True
    close[ceiling_251,ceiling_58]=True
    close[ceiling_251,wall_69]=True
    close[ceiling_251,wall_244]=True
    close[ceiling_251,wall_246]=True
    close[ceiling_251,wall_247]=True
    close[ceiling_251,ceiling_250]=True
    close[ceiling_251,ceiling_252]=True
    close[ceiling_251,ceiling_254]=True
    close[ceiling_251,light_283]=True
    close[ceiling_251,ceilinglamp_303]=True
    close[ceiling_251,doorjamb_309]=True
    close[ceiling_252,ceiling_59]=True
    close[ceiling_252,wall_65]=True
    close[ceiling_252,wall_246]=True
    close[ceiling_252,ceiling_251]=True
    close[ceiling_252,ceiling_253]=True
    close[ceiling_252,chair_271]=True
    close[ceiling_252,bookshelf_275]=True
    close[ceiling_252,cpuscreen_277]=True
    close[ceiling_252,walllamp_304]=True
    close[ceiling_253,wall_243]=True
    close[ceiling_253,wall_246]=True
    close[ceiling_253,wall_249]=True
    close[ceiling_253,ceiling_252]=True
    close[ceiling_253,ceiling_254]=True
    close[ceiling_253,ceiling_258]=True
    close[ceiling_253,chair_271]=True
    close[ceiling_253,cpuscreen_277]=True
    close[ceiling_253,ceilinglamp_303]=True
    close[ceiling_253,walllamp_304]=True
    close[ceiling_253,walllamp_305]=True
    close[ceiling_254,ceiling_251]=True
    close[ceiling_254,ceiling_253]=True
    close[ceiling_254,ceiling_255]=True
    close[ceiling_254,ceiling_257]=True
    close[ceiling_254,ceilinglamp_303]=True
    close[ceiling_255,wall_242]=True
    close[ceiling_255,wall_247]=True
    close[ceiling_255,wall_248]=True
    close[ceiling_255,ceiling_250]=True
    close[ceiling_255,ceiling_254]=True
    close[ceiling_255,ceiling_256]=True
    close[ceiling_255,drawing_288]=True
    close[ceiling_255,ceilinglamp_303]=True
    close[ceiling_255,walllamp_306]=True
    close[ceiling_255,walllamp_307]=True
    close[ceiling_256,wall_248]=True
    close[ceiling_256,ceiling_255]=True
    close[ceiling_256,ceiling_257]=True
    close[ceiling_256,curtain_291]=True
    close[ceiling_256,walllamp_307]=True
    close[ceiling_257,wall_245]=True
    close[ceiling_257,wall_248]=True
    close[ceiling_257,wall_249]=True
    close[ceiling_257,ceiling_254]=True
    close[ceiling_257,ceiling_256]=True
    close[ceiling_257,ceiling_258]=True
    close[ceiling_257,curtain_289]=True
    close[ceiling_257,curtain_290]=True
    close[ceiling_257,curtain_291]=True
    close[ceiling_257,hanger_292]=True
    close[ceiling_257,hanger_293]=True
    close[ceiling_257,hanger_294]=True
    close[ceiling_257,ceilinglamp_303]=True
    close[ceiling_257,window_310]=True
    close[ceiling_258,wall_249]=True
    close[ceiling_258,ceiling_253]=True
    close[ceiling_258,ceiling_257]=True
    close[ceiling_258,dresser_274]=True
    close[ceiling_258,curtain_289]=True
    close[ceiling_258,curtain_290]=True
    close[ceiling_258,hanger_292]=True
    close[ceiling_258,hanger_293]=True
    close[ceiling_258,hanger_294]=True
    close[ceiling_258,walllamp_305]=True
    close[ceiling_258,doorjamb_308]=True
    close[floor_259,door_62]=True
    close[floor_259,wall_247]=True
    close[floor_259,floor_260]=True
    close[floor_259,floor_261]=True
    close[floor_259,floor_265]=True
    close[floor_259,tvstand_273]=True
    close[floor_259,television_281]=True
    close[floor_259,powersocket_282]=True
    close[floor_259,mat_284]=True
    close[floor_259,walllamp_306]=True
    close[floor_260,door_62]=True
    close[floor_260,wall_247]=True
    close[floor_260,floor_259]=True
    close[floor_260,floor_261]=True
    close[floor_260,floor_265]=True
    close[floor_260,tvstand_273]=True
    close[floor_260,television_281]=True
    close[floor_260,powersocket_282]=True
    close[floor_260,mat_284]=True
    close[floor_260,walllamp_306]=True
    close[floor_261,floor_49]=True
    close[floor_261,door_62]=True
    close[floor_261,wall_69]=True
    close[floor_261,wall_244]=True
    close[floor_261,wall_246]=True
    close[floor_261,wall_247]=True
    close[floor_261,floor_259]=True
    close[floor_261,floor_260]=True
    close[floor_261,floor_262]=True
    close[floor_261,floor_264]=True
    close[floor_261,chair_271]=True
    close[floor_261,tvstand_273]=True
    close[floor_261,television_281]=True
    close[floor_261,powersocket_282]=True
    close[floor_261,light_283]=True
    close[floor_261,mat_284]=True
    close[floor_261,doorjamb_309]=True
    close[floor_262,floor_50]=True
    close[floor_262,door_62]=True
    close[floor_262,wall_65]=True
    close[floor_262,trashcan_99]=True
    close[floor_262,wall_246]=True
    close[floor_262,floor_261]=True
    close[floor_262,floor_263]=True
    close[floor_262,chair_271]=True
    close[floor_262,desk_272]=True
    close[floor_262,bookshelf_275]=True
    close[floor_262,computer_276]=True
    close[floor_262,cpuscreen_277]=True
    close[floor_262,keyboard_278]=True
    close[floor_262,light_283]=True
    close[floor_262,mat_284]=True
    close[floor_262,walllamp_304]=True
    close[floor_263,wall_243]=True
    close[floor_263,wall_246]=True
    close[floor_263,wall_249]=True
    close[floor_263,floor_262]=True
    close[floor_263,floor_264]=True
    close[floor_263,floor_268]=True
    close[floor_263,chair_271]=True
    close[floor_263,desk_272]=True
    close[floor_263,computer_276]=True
    close[floor_263,cpuscreen_277]=True
    close[floor_263,keyboard_278]=True
    close[floor_263,mousepad_279]=True
    close[floor_263,mouse_280]=True
    close[floor_263,walllamp_305]=True
    close[floor_264,floor_261]=True
    close[floor_264,floor_263]=True
    close[floor_264,floor_265]=True
    close[floor_264,floor_267]=True
    close[floor_264,couch_269]=True
    close[floor_264,table_270]=True
    close[floor_264,chair_271]=True
    close[floor_264,mat_284]=True
    close[floor_264,orchid_285]=True
    close[floor_265,wall_242]=True
    close[floor_265,wall_247]=True
    close[floor_265,wall_248]=True
    close[floor_265,floor_259]=True
    close[floor_265,floor_260]=True
    close[floor_265,floor_264]=True
    close[floor_265,floor_266]=True
    close[floor_265,couch_269]=True
    close[floor_265,table_270]=True
    close[floor_265,orchid_285]=True
    close[floor_265,drawing_288]=True
    close[floor_265,walllamp_307]=True
    close[floor_266,wall_248]=True
    close[floor_266,floor_265]=True
    close[floor_266,floor_267]=True
    close[floor_266,couch_269]=True
    close[floor_266,table_270]=True
    close[floor_266,orchid_285]=True
    close[floor_266,pillow_286]=True
    close[floor_266,pillow_287]=True
    close[floor_267,wall_245]=True
    close[floor_267,wall_248]=True
    close[floor_267,wall_249]=True
    close[floor_267,floor_264]=True
    close[floor_267,floor_266]=True
    close[floor_267,floor_268]=True
    close[floor_267,couch_269]=True
    close[floor_267,table_270]=True
    close[floor_267,dresser_274]=True
    close[floor_267,orchid_285]=True
    close[floor_267,pillow_286]=True
    close[floor_267,pillow_287]=True
    close[floor_267,curtain_289]=True
    close[floor_267,curtain_290]=True
    close[floor_267,curtain_291]=True
    close[floor_267,window_310]=True
    close[floor_268,wall_249]=True
    close[floor_268,floor_263]=True
    close[floor_268,floor_267]=True
    close[floor_268,dresser_274]=True
    close[floor_268,computer_276]=True
    close[floor_268,doorjamb_308]=True
    close[couch_269,wall_242]=True
    close[couch_269,wall_245]=True
    close[couch_269,wall_248]=True
    close[couch_269,floor_264]=True
    close[couch_269,floor_265]=True
    close[couch_269,floor_266]=True
    close[couch_269,floor_267]=True
    close[couch_269,table_270]=True
    close[couch_269,orchid_285]=True
    close[couch_269,pillow_286]=True
    close[couch_269,pillow_287]=True
    close[couch_269,drawing_288]=True
    close[couch_269,curtain_289]=True
    close[couch_269,curtain_290]=True
    close[couch_269,curtain_291]=True
    close[couch_269,ceilinglamp_303]=True
    close[couch_269,walllamp_307]=True
    close[couch_269,window_310]=True
    close[couch_269,brush_2002]=True
    close[couch_269,phone_2017]=True
    close[couch_269,shoes_2033]=True
    close[table_270,wall_248]=True
    close[table_270,floor_264]=True
    close[table_270,floor_265]=True
    close[table_270,floor_266]=True
    close[table_270,floor_267]=True
    close[table_270,couch_269]=True
    close[table_270,orchid_285]=True
    close[table_270,pillow_286]=True
    close[table_270,pillow_287]=True
    close[table_270,pencil_2014]=True
    close[table_270,shampoo_2019]=True
    close[chair_271,wall_246]=True
    close[chair_271,ceiling_252]=True
    close[chair_271,ceiling_253]=True
    close[chair_271,floor_261]=True
    close[chair_271,floor_262]=True
    close[chair_271,floor_263]=True
    close[chair_271,floor_264]=True
    close[chair_271,desk_272]=True
    close[chair_271,computer_276]=True
    close[chair_271,cpuscreen_277]=True
    close[chair_271,keyboard_278]=True
    close[chair_271,mousepad_279]=True
    close[chair_271,mouse_280]=True
    close[chair_271,mat_284]=True
    close[chair_271,walllamp_304]=True
    close[desk_272,headset_2146]=True
    close[desk_272,phone_2147]=True
    close[desk_272,wall_243]=True
    close[desk_272,wall_246]=True
    close[desk_272,floor_262]=True
    close[desk_272,floor_263]=True
    close[desk_272,chair_271]=True
    close[desk_272,computer_276]=True
    close[desk_272,cpuscreen_277]=True
    close[desk_272,keyboard_278]=True
    close[desk_272,mousepad_279]=True
    close[desk_272,mouse_280]=True
    close[desk_272,walllamp_304]=True
    close[desk_272,walllamp_305]=True
    close[desk_272,stamp_2022]=True
    close[desk_272,stamp_2043]=True
    close[tvstand_273,remote_control_2124]=True
    close[tvstand_273,cd_player_2129]=True
    close[tvstand_273,dvd_player_2130]=True
    close[tvstand_273,headset_2131]=True
    close[tvstand_273,cd_2145]=True
    close[tvstand_273,floor_49]=True
    close[tvstand_273,door_62]=True
    close[tvstand_273,wall_69]=True
    close[tvstand_273,wall_244]=True
    close[tvstand_273,wall_247]=True
    close[tvstand_273,floor_259]=True
    close[tvstand_273,floor_260]=True
    close[tvstand_273,floor_261]=True
    close[tvstand_273,television_281]=True
    close[tvstand_273,powersocket_282]=True
    close[tvstand_273,mat_284]=True
    close[tvstand_273,doorjamb_309]=True
    close[dresser_274,wall_245]=True
    close[dresser_274,wall_249]=True
    close[dresser_274,ceiling_258]=True
    close[dresser_274,floor_267]=True
    close[dresser_274,floor_268]=True
    close[dresser_274,curtain_289]=True
    close[dresser_274,curtain_290]=True
    close[dresser_274,hanger_292]=True
    close[dresser_274,hanger_293]=True
    close[dresser_274,hanger_294]=True
    close[dresser_274,doorjamb_308]=True
    close[dresser_274,window_310]=True
    close[dresser_274,blow_dryer_2057]=True
    close[dresser_274,cat_2069]=True
    close[dresser_274,check_2075]=True
    close[bookshelf_275,floor_50]=True
    close[bookshelf_275,floor_51]=True
    close[bookshelf_275,ceiling_59]=True
    close[bookshelf_275,wall_65]=True
    close[bookshelf_275,wall_68]=True
    close[bookshelf_275,trashcan_99]=True
    close[bookshelf_275,wall_246]=True
    close[bookshelf_275,ceiling_252]=True
    close[bookshelf_275,floor_262]=True
    close[bookshelf_275,pencil_2020]=True
    close[computer_276,wall_243]=True
    close[computer_276,wall_246]=True
    close[computer_276,wall_249]=True
    close[computer_276,floor_262]=True
    close[computer_276,floor_263]=True
    close[computer_276,floor_268]=True
    close[computer_276,chair_271]=True
    close[computer_276,desk_272]=True
    close[computer_276,cpuscreen_277]=True
    close[computer_276,keyboard_278]=True
    close[computer_276,mousepad_279]=True
    close[computer_276,mouse_280]=True
    close[computer_276,walllamp_305]=True
    close[cpuscreen_277,wall_243]=True
    close[cpuscreen_277,wall_246]=True
    close[cpuscreen_277,ceiling_252]=True
    close[cpuscreen_277,ceiling_253]=True
    close[cpuscreen_277,floor_262]=True
    close[cpuscreen_277,floor_263]=True
    close[cpuscreen_277,chair_271]=True
    close[cpuscreen_277,desk_272]=True
    close[cpuscreen_277,computer_276]=True
    close[cpuscreen_277,keyboard_278]=True
    close[cpuscreen_277,mousepad_279]=True
    close[cpuscreen_277,mouse_280]=True
    close[cpuscreen_277,walllamp_304]=True
    close[cpuscreen_277,walllamp_305]=True
    close[keyboard_278,wall_243]=True
    close[keyboard_278,wall_246]=True
    close[keyboard_278,floor_262]=True
    close[keyboard_278,floor_263]=True
    close[keyboard_278,chair_271]=True
    close[keyboard_278,desk_272]=True
    close[keyboard_278,computer_276]=True
    close[keyboard_278,cpuscreen_277]=True
    close[keyboard_278,mousepad_279]=True
    close[keyboard_278,mouse_280]=True
    close[keyboard_278,walllamp_304]=True
    close[keyboard_278,walllamp_305]=True
    close[mousepad_279,wall_243]=True
    close[mousepad_279,wall_246]=True
    close[mousepad_279,wall_249]=True
    close[mousepad_279,floor_263]=True
    close[mousepad_279,chair_271]=True
    close[mousepad_279,desk_272]=True
    close[mousepad_279,computer_276]=True
    close[mousepad_279,cpuscreen_277]=True
    close[mousepad_279,keyboard_278]=True
    close[mousepad_279,mouse_280]=True
    close[mousepad_279,walllamp_305]=True
    close[mouse_280,wall_243]=True
    close[mouse_280,wall_246]=True
    close[mouse_280,wall_249]=True
    close[mouse_280,floor_263]=True
    close[mouse_280,chair_271]=True
    close[mouse_280,desk_272]=True
    close[mouse_280,computer_276]=True
    close[mouse_280,cpuscreen_277]=True
    close[mouse_280,keyboard_278]=True
    close[mouse_280,mousepad_279]=True
    close[mouse_280,walllamp_305]=True
    close[television_281,door_62]=True
    close[television_281,wall_69]=True
    close[television_281,wall_244]=True
    close[television_281,wall_247]=True
    close[television_281,ceiling_250]=True
    close[television_281,floor_259]=True
    close[television_281,floor_260]=True
    close[television_281,floor_261]=True
    close[television_281,tvstand_273]=True
    close[television_281,powersocket_282]=True
    close[television_281,doorjamb_309]=True
    close[powersocket_282,floor_49]=True
    close[powersocket_282,door_62]=True
    close[powersocket_282,wall_69]=True
    close[powersocket_282,wall_244]=True
    close[powersocket_282,wall_247]=True
    close[powersocket_282,floor_259]=True
    close[powersocket_282,floor_260]=True
    close[powersocket_282,floor_261]=True
    close[powersocket_282,tvstand_273]=True
    close[powersocket_282,television_281]=True
    close[powersocket_282,light_283]=True
    close[powersocket_282,mat_284]=True
    close[powersocket_282,doorjamb_309]=True
    close[light_283,floor_49]=True
    close[light_283,floor_50]=True
    close[light_283,ceiling_58]=True
    close[light_283,door_62]=True
    close[light_283,wall_65]=True
    close[light_283,wall_69]=True
    close[light_283,wall_244]=True
    close[light_283,wall_246]=True
    close[light_283,ceiling_251]=True
    close[light_283,floor_261]=True
    close[light_283,floor_262]=True
    close[light_283,powersocket_282]=True
    close[light_283,mat_284]=True
    close[light_283,doorjamb_309]=True
    close[mat_284,floor_49]=True
    close[mat_284,door_62]=True
    close[mat_284,wall_69]=True
    close[mat_284,wall_244]=True
    close[mat_284,wall_246]=True
    close[mat_284,wall_247]=True
    close[mat_284,floor_259]=True
    close[mat_284,floor_260]=True
    close[mat_284,floor_261]=True
    close[mat_284,floor_262]=True
    close[mat_284,floor_264]=True
    close[mat_284,chair_271]=True
    close[mat_284,tvstand_273]=True
    close[mat_284,powersocket_282]=True
    close[mat_284,light_283]=True
    close[mat_284,doorjamb_309]=True
    close[orchid_285,wall_248]=True
    close[orchid_285,floor_264]=True
    close[orchid_285,floor_265]=True
    close[orchid_285,floor_266]=True
    close[orchid_285,floor_267]=True
    close[orchid_285,couch_269]=True
    close[orchid_285,table_270]=True
    close[orchid_285,pillow_287]=True
    close[pillow_286,wall_245]=True
    close[pillow_286,wall_248]=True
    close[pillow_286,floor_266]=True
    close[pillow_286,floor_267]=True
    close[pillow_286,couch_269]=True
    close[pillow_286,table_270]=True
    close[pillow_286,pillow_287]=True
    close[pillow_286,curtain_291]=True
    close[pillow_286,window_310]=True
    close[pillow_287,wall_245]=True
    close[pillow_287,wall_248]=True
    close[pillow_287,floor_266]=True
    close[pillow_287,floor_267]=True
    close[pillow_287,couch_269]=True
    close[pillow_287,table_270]=True
    close[pillow_287,orchid_285]=True
    close[pillow_287,pillow_286]=True
    close[pillow_287,curtain_289]=True
    close[pillow_287,curtain_290]=True
    close[pillow_287,curtain_291]=True
    close[pillow_287,window_310]=True
    close[drawing_288,wall_242]=True
    close[drawing_288,wall_247]=True
    close[drawing_288,ceiling_250]=True
    close[drawing_288,ceiling_255]=True
    close[drawing_288,floor_265]=True
    close[drawing_288,couch_269]=True
    close[drawing_288,walllamp_306]=True
    close[drawing_288,walllamp_307]=True
    close[curtain_289,wall_245]=True
    close[curtain_289,wall_249]=True
    close[curtain_289,ceiling_257]=True
    close[curtain_289,ceiling_258]=True
    close[curtain_289,floor_267]=True
    close[curtain_289,couch_269]=True
    close[curtain_289,dresser_274]=True
    close[curtain_289,pillow_287]=True
    close[curtain_289,curtain_290]=True
    close[curtain_289,curtain_291]=True
    close[curtain_289,hanger_292]=True
    close[curtain_289,hanger_293]=True
    close[curtain_289,hanger_294]=True
    close[curtain_289,window_310]=True
    close[curtain_290,wall_245]=True
    close[curtain_290,wall_249]=True
    close[curtain_290,ceiling_257]=True
    close[curtain_290,ceiling_258]=True
    close[curtain_290,floor_267]=True
    close[curtain_290,couch_269]=True
    close[curtain_290,dresser_274]=True
    close[curtain_290,pillow_287]=True
    close[curtain_290,curtain_289]=True
    close[curtain_290,curtain_291]=True
    close[curtain_290,hanger_292]=True
    close[curtain_290,hanger_293]=True
    close[curtain_290,hanger_294]=True
    close[curtain_290,window_310]=True
    close[curtain_291,wall_245]=True
    close[curtain_291,wall_248]=True
    close[curtain_291,ceiling_256]=True
    close[curtain_291,ceiling_257]=True
    close[curtain_291,floor_267]=True
    close[curtain_291,couch_269]=True
    close[curtain_291,pillow_286]=True
    close[curtain_291,pillow_287]=True
    close[curtain_291,curtain_289]=True
    close[curtain_291,curtain_290]=True
    close[curtain_291,window_310]=True
    close[hanger_292,wall_245]=True
    close[hanger_292,wall_249]=True
    close[hanger_292,ceiling_257]=True
    close[hanger_292,ceiling_258]=True
    close[hanger_292,dresser_274]=True
    close[hanger_292,curtain_289]=True
    close[hanger_292,curtain_290]=True
    close[hanger_292,hanger_293]=True
    close[hanger_292,hanger_294]=True
    close[hanger_292,window_310]=True
    close[hanger_292,clothes_pants_2036]=True
    close[hanger_293,wall_245]=True
    close[hanger_293,wall_249]=True
    close[hanger_293,ceiling_257]=True
    close[hanger_293,ceiling_258]=True
    close[hanger_293,dresser_274]=True
    close[hanger_293,curtain_289]=True
    close[hanger_293,curtain_290]=True
    close[hanger_293,hanger_292]=True
    close[hanger_293,hanger_294]=True
    close[hanger_293,window_310]=True
    close[hanger_294,wall_245]=True
    close[hanger_294,wall_249]=True
    close[hanger_294,ceiling_257]=True
    close[hanger_294,ceiling_258]=True
    close[hanger_294,dresser_274]=True
    close[hanger_294,curtain_289]=True
    close[hanger_294,curtain_290]=True
    close[hanger_294,hanger_292]=True
    close[hanger_294,hanger_293]=True
    close[hanger_294,window_310]=True
    close[ceilinglamp_303,ceiling_251]=True
    close[ceilinglamp_303,ceiling_253]=True
    close[ceilinglamp_303,ceiling_254]=True
    close[ceilinglamp_303,ceiling_255]=True
    close[ceilinglamp_303,ceiling_257]=True
    close[ceilinglamp_303,couch_269]=True
    close[walllamp_304,wall_243]=True
    close[walllamp_304,wall_246]=True
    close[walllamp_304,ceiling_252]=True
    close[walllamp_304,ceiling_253]=True
    close[walllamp_304,floor_262]=True
    close[walllamp_304,chair_271]=True
    close[walllamp_304,desk_272]=True
    close[walllamp_304,cpuscreen_277]=True
    close[walllamp_304,keyboard_278]=True
    close[walllamp_305,wall_243]=True
    close[walllamp_305,wall_249]=True
    close[walllamp_305,ceiling_253]=True
    close[walllamp_305,ceiling_258]=True
    close[walllamp_305,floor_263]=True
    close[walllamp_305,desk_272]=True
    close[walllamp_305,computer_276]=True
    close[walllamp_305,cpuscreen_277]=True
    close[walllamp_305,keyboard_278]=True
    close[walllamp_305,mousepad_279]=True
    close[walllamp_305,mouse_280]=True
    close[walllamp_306,wall_242]=True
    close[walllamp_306,wall_247]=True
    close[walllamp_306,ceiling_250]=True
    close[walllamp_306,ceiling_255]=True
    close[walllamp_306,floor_259]=True
    close[walllamp_306,floor_260]=True
    close[walllamp_306,drawing_288]=True
    close[walllamp_307,wall_242]=True
    close[walllamp_307,wall_248]=True
    close[walllamp_307,ceiling_255]=True
    close[walllamp_307,ceiling_256]=True
    close[walllamp_307,floor_265]=True
    close[walllamp_307,couch_269]=True
    close[walllamp_307,drawing_288]=True
    close[doorjamb_308,wall_243]=True
    close[doorjamb_308,wall_249]=True
    close[doorjamb_308,ceiling_258]=True
    close[doorjamb_308,floor_268]=True
    close[doorjamb_308,dresser_274]=True
    close[doorjamb_309,floor_49]=True
    close[doorjamb_309,ceiling_58]=True
    close[doorjamb_309,door_62]=True
    close[doorjamb_309,wall_65]=True
    close[doorjamb_309,wall_69]=True
    close[doorjamb_309,wall_244]=True
    close[doorjamb_309,wall_246]=True
    close[doorjamb_309,wall_247]=True
    close[doorjamb_309,ceiling_251]=True
    close[doorjamb_309,floor_261]=True
    close[doorjamb_309,tvstand_273]=True
    close[doorjamb_309,television_281]=True
    close[doorjamb_309,powersocket_282]=True
    close[doorjamb_309,light_283]=True
    close[doorjamb_309,mat_284]=True
    close[window_310,wall_245]=True
    close[window_310,wall_248]=True
    close[window_310,wall_249]=True
    close[window_310,ceiling_257]=True
    close[window_310,floor_267]=True
    close[window_310,couch_269]=True
    close[window_310,dresser_274]=True
    close[window_310,pillow_286]=True
    close[window_310,pillow_287]=True
    close[window_310,curtain_289]=True
    close[window_310,curtain_290]=True
    close[window_310,curtain_291]=True
    close[window_310,hanger_292]=True
    close[window_310,hanger_293]=True
    close[window_310,hanger_294]=True
    close[food_food_1000,fridge_126]=True
    close[wooden_spoon_2000,table_199]=True
    close[food_food_2001,fridge_126]=True
    close[brush_2002,couch_269]=True
    close[chair_2003,couch_198]=True
    close[lighter_2004,mat_102]=True
    close[table_cloth_2005,table_114]=True
    close[table_cloth_2005,food_butter_2007]=True
    close[piano_bench_2006,floor_44]=True
    close[food_butter_2007,table_cloth_2005]=True
    close[diary_2008,filing_cabinet_200]=True
    close[food_onion_2009,trashcan_99]=True
    close[soap_2010,sink_120]=True
    close[detergent_2011,dishwasher_129]=True
    close[measuring_cup_2012,dishwasher_129]=True
    close[oil_2013,oven_127]=True
    close[pencil_2014,table_270]=True
    close[food_carrot_2015,oven_127]=True
    close[phone_2016,couch_198]=True
    close[phone_2017,couch_269]=True
    close[envelope_2018,filing_cabinet_200]=True
    close[shampoo_2019,table_270]=True
    close[pencil_2020,bookshelf_275]=True
    close[food_food_2021,table_114]=True
    close[stamp_2022,desk_272]=True
    close[tea_bag_2023,table_199]=True
    close[ice_2024,sink_120]=True
    close[rag_2025,filing_cabinet_200]=True
    close[check_2026,desk_193]=True
    close[food_orange_2027,kitchen_counter_123]=True
    close[instrument_guitar_2028,couch_198]=True
    close[phone_2029,bathroom_counter_18]=True
    close[cd_2030,filing_cabinet_200]=True
    close[scrabble_2031,filing_cabinet_200]=True
    close[shoes_2033,couch_269]=True
    close[laser_pointer_2034,desk_193]=True
    close[knife_2035,kitchen_counter_123]=True
    close[clothes_pants_2036,hanger_292]=True
    close[knife_2037,cupboard_118]=True
    close[box_2038,table_114]=True
    close[lighter_2039,mat_102]=True
    close[pot_2040,microwave_135]=True
    close[food_salt_2041,kitchen_counter_119]=True
    close[after_shave_2042,filing_cabinet_200]=True
    close[stamp_2043,desk_272]=True
    close[shoe_rack_2044,mat_203]=True
    close[shoe_rack_2044,chessboard_2070]=True
    close[shoe_rack_2044,check_2071]=True
    close[glue_2045,trashcan_99]=True
    close[food_food_2046,fridge_126]=True
    close[homework_2047,filing_cabinet_200]=True
    close[food_onion_2048,fridge_126]=True
    close[cup_2049,table_114]=True
    close[stereo_2050,filing_cabinet_200]=True
    close[after_shave_2051,filing_cabinet_200]=True
    close[rag_2052,couch_198]=True
    close[coffee_filter_2053,cupboard_117]=True
    close[food_kiwi_2054,kitchen_counter_123]=True
    close[envelope_2055,bookshelf_124]=True
    close[toy_2056,mat_32]=True
    close[blow_dryer_2057,dresser_274]=True
    close[check_2058,table_114]=True
    close[tooth_paste_2059,bathroom_cabinet_17]=True
    close[novel_2060,bookshelf_196]=True
    close[food_orange_2061,trashcan_99]=True
    close[piano_bench_2062,floor_44]=True
    close[after_shave_2063,sink_19]=True
    close[food_food_2064,oven_127]=True
    close[coffee_filter_2065,coffe_maker_130]=True
    close[tea_2066,cupboard_118]=True
    close[piano_bench_2067,mat_32]=True
    close[tray_2068,kitchen_counter_123]=True
    close[cat_2069,dresser_274]=True
    close[chessboard_2070,shoe_rack_2044]=True
    close[check_2071,shoe_rack_2044]=True
    close[food_cheese_2072,oven_127]=True
    close[food_food_2073,fridge_126]=True
    close[food_food_2074,filing_cabinet_200]=True
    close[check_2075,dresser_274]=True
    close[toilet_paper_2076,toilet_15]=True
    close[food_peanut_butter_2077,cupboard_118]=True
    facing[wall_2,drawing_33]=True
    facing[wall_2,drawing_110]=True
    facing[wall_3,drawing_33]=True
    facing[wall_4,drawing_33]=True
    facing[wall_5,drawing_33]=True
    facing[ceiling_6,drawing_33]=True
    facing[ceiling_7,drawing_33]=True
    facing[ceiling_7,drawing_110]=True
    facing[ceiling_8,drawing_33]=True
    facing[ceiling_9,drawing_33]=True
    facing[floor_10,drawing_33]=True
    facing[floor_11,drawing_33]=True
    facing[floor_12,drawing_33]=True
    facing[floor_12,drawing_110]=True
    facing[floor_13,drawing_33]=True
    facing[floor_14,drawing_33]=True
    facing[toilet_15,drawing_33]=True
    facing[shower_16,drawing_33]=True
    facing[bathroom_cabinet_17,drawing_33]=True
    facing[bathroom_counter_18,drawing_33]=True
    facing[sink_19,drawing_33]=True
    facing[faucet_20,drawing_33]=True
    facing[shower_21,drawing_33]=True
    facing[curtain_22,drawing_33]=True
    facing[mat_32,drawing_33]=True
    facing[walllamp_34,drawing_33]=True
    facing[ceilinglamp_35,drawing_33]=True
    facing[walllamp_36,drawing_33]=True
    facing[doorjamb_37,drawing_110]=True
    facing[door_38,drawing_110]=True
    facing[floor_42,drawing_110]=True
    facing[floor_42,drawing_111]=True
    facing[floor_43,drawing_110]=True
    facing[floor_43,drawing_111]=True
    facing[floor_44,drawing_110]=True
    facing[floor_44,drawing_111]=True
    facing[floor_47,drawing_110]=True
    facing[floor_47,drawing_111]=True
    facing[floor_48,drawing_110]=True
    facing[floor_48,drawing_111]=True
    facing[floor_49,drawing_111]=True
    facing[floor_50,drawing_111]=True
    facing[ceiling_52,drawing_110]=True
    facing[ceiling_52,drawing_111]=True
    facing[ceiling_53,drawing_110]=True
    facing[ceiling_53,drawing_111]=True
    facing[ceiling_56,drawing_110]=True
    facing[ceiling_56,drawing_111]=True
    facing[ceiling_57,drawing_110]=True
    facing[ceiling_57,drawing_111]=True
    facing[ceiling_58,drawing_111]=True
    facing[ceiling_59,drawing_111]=True
    facing[door_61,drawing_202]=True
    facing[door_62,drawing_111]=True
    facing[door_62,computer_276]=True
    facing[door_62,drawing_288]=True
    facing[wall_63,drawing_110]=True
    facing[wall_66,drawing_202]=True
    facing[wall_69,drawing_111]=True
    facing[wall_70,drawing_110]=True
    facing[wall_70,drawing_111]=True
    facing[mat_102,drawing_110]=True
    facing[mat_102,drawing_111]=True
    facing[pillow_103,drawing_110]=True
    facing[pillow_103,drawing_111]=True
    facing[pillow_104,drawing_110]=True
    facing[pillow_104,drawing_111]=True
    facing[pillow_105,drawing_110]=True
    facing[pillow_105,drawing_111]=True
    facing[pillow_106,drawing_110]=True
    facing[pillow_106,drawing_111]=True
    facing[pillow_107,drawing_110]=True
    facing[pillow_107,drawing_111]=True
    facing[pillow_108,drawing_110]=True
    facing[pillow_108,drawing_111]=True
    facing[drawing_110,drawing_111]=True
    facing[drawing_111,drawing_110]=True
    facing[bench_113,drawing_110]=True
    facing[table_114,drawing_110]=True
    facing[table_114,drawing_111]=True
    facing[bench_115,drawing_110]=True
    facing[bench_115,drawing_111]=True
    facing[tvstand_116,drawing_110]=True
    facing[tvstand_116,drawing_111]=True
    facing[bookshelf_124,drawing_110]=True
    facing[bookshelf_124,drawing_111]=True
    facing[ceilinglamp_137,drawing_110]=True
    facing[ceilinglamp_137,drawing_111]=True
    facing[ceilinglamp_138,drawing_111]=True
    facing[floor_163,drawing_201]=True
    facing[floor_163,computer_209]=True
    facing[floor_164,drawing_201]=True
    facing[floor_164,computer_209]=True
    facing[floor_165,drawing_201]=True
    facing[floor_165,computer_209]=True
    facing[floor_166,drawing_201]=True
    facing[floor_167,drawing_201]=True
    facing[floor_168,drawing_201]=True
    facing[floor_168,drawing_202]=True
    facing[floor_168,computer_209]=True
    facing[floor_169,drawing_202]=True
    facing[floor_169,computer_209]=True
    facing[floor_170,drawing_202]=True
    facing[floor_171,drawing_202]=True
    facing[floor_171,computer_209]=True
    facing[floor_172,drawing_202]=True
    facing[wall_173,computer_209]=True
    facing[wall_175,drawing_201]=True
    facing[wall_175,computer_209]=True
    facing[wall_176,drawing_202]=True
    facing[wall_177,drawing_202]=True
    facing[wall_178,drawing_201]=True
    facing[wall_179,drawing_202]=True
    facing[wall_180,drawing_201]=True
    facing[ceiling_181,computer_209]=True
    facing[ceiling_182,drawing_202]=True
    facing[ceiling_182,computer_209]=True
    facing[ceiling_183,drawing_202]=True
    facing[ceiling_184,drawing_202]=True
    facing[ceiling_185,drawing_201]=True
    facing[ceiling_185,drawing_202]=True
    facing[ceiling_185,computer_209]=True
    facing[ceiling_186,drawing_201]=True
    facing[ceiling_186,computer_209]=True
    facing[ceiling_187,drawing_201]=True
    facing[ceiling_188,drawing_201]=True
    facing[ceiling_189,drawing_202]=True
    facing[doorjamb_190,drawing_202]=True
    facing[window_191,drawing_201]=True
    facing[nightstand_192,drawing_201]=True
    facing[chair_194,computer_209]=True
    facing[nightstand_195,drawing_201]=True
    facing[nightstand_195,computer_209]=True
    facing[bookshelf_196,drawing_202]=True
    facing[bed_197,computer_209]=True
    facing[table_199,drawing_201]=True
    facing[table_199,drawing_202]=True
    facing[table_199,computer_209]=True
    facing[filing_cabinet_200,drawing_202]=True
    facing[mat_203,drawing_202]=True
    facing[curtain_204,drawing_201]=True
    facing[curtain_205,drawing_201]=True
    facing[curtain_206,drawing_201]=True
    facing[pillow_207,drawing_201]=True
    facing[pillow_208,drawing_201]=True
    facing[keyboard_211,drawing_201]=True
    facing[light_212,drawing_202]=True
    facing[photoframe_219,drawing_202]=True
    facing[ceilinglamp_237,drawing_201]=True
    facing[ceilinglamp_237,drawing_202]=True
    facing[tablelamp_238,drawing_201]=True
    facing[tablelamp_239,drawing_201]=True
    facing[tablelamp_239,computer_209]=True
    facing[wall_242,television_281]=True
    facing[wall_244,drawing_111]=True
    facing[wall_244,drawing_288]=True
    facing[wall_245,computer_276]=True
    facing[wall_247,television_281]=True
    facing[wall_247,drawing_288]=True
    facing[wall_248,drawing_288]=True
    facing[ceiling_250,television_281]=True
    facing[ceiling_250,drawing_288]=True
    facing[ceiling_251,computer_276]=True
    facing[ceiling_251,television_281]=True
    facing[ceiling_251,drawing_288]=True
    facing[ceiling_253,computer_276]=True
    facing[ceiling_254,computer_276]=True
    facing[ceiling_254,television_281]=True
    facing[ceiling_254,drawing_288]=True
    facing[ceiling_255,television_281]=True
    facing[ceiling_255,drawing_288]=True
    facing[ceiling_256,drawing_288]=True
    facing[ceiling_257,computer_276]=True
    facing[ceiling_257,drawing_288]=True
    facing[floor_259,television_281]=True
    facing[floor_259,drawing_288]=True
    facing[floor_260,television_281]=True
    facing[floor_260,drawing_288]=True
    facing[floor_261,computer_276]=True
    facing[floor_261,television_281]=True
    facing[floor_261,drawing_288]=True
    facing[floor_263,computer_276]=True
    facing[floor_264,computer_276]=True
    facing[floor_264,television_281]=True
    facing[floor_264,drawing_288]=True
    facing[floor_265,television_281]=True
    facing[floor_265,drawing_288]=True
    facing[floor_267,computer_276]=True
    facing[floor_267,drawing_288]=True
    facing[couch_269,drawing_288]=True
    facing[table_270,computer_276]=True
    facing[table_270,television_281]=True
    facing[table_270,drawing_288]=True
    facing[chair_271,computer_276]=True
    facing[tvstand_273,television_281]=True
    facing[tvstand_273,drawing_288]=True
    facing[mousepad_279,computer_276]=True
    facing[television_281,drawing_288]=True
    facing[mat_284,computer_276]=True
    facing[mat_284,television_281]=True
    facing[mat_284,drawing_288]=True
    facing[orchid_285,computer_276]=True
    facing[orchid_285,television_281]=True
    facing[orchid_285,drawing_288]=True
    facing[pillow_286,drawing_288]=True
    facing[pillow_287,drawing_288]=True
    facing[drawing_288,television_281]=True
    facing[ceilinglamp_303,computer_276]=True
    facing[ceilinglamp_303,television_281]=True
    facing[ceilinglamp_303,drawing_288]=True
    facing[walllamp_306,television_281]=True
    facing[walllamp_307,television_281]=True
    facing[doorjamb_309,drawing_111]=True
    facing[doorjamb_309,drawing_288]=True
    #relations_end

    #exploration
    #exploration_end

    #id
    id[clothes_pants_2157]=2157
    id[clothes_shirt_2158]=2158
    id[clothes_socks_2159]=2159
    id[clothes_skirt_2160]=2160
    id[iron_2161]=2161
    id[basket_for_clothes_2078]=2078
    id[washing_machine_2079]=2079
    id[food_steak_2080]=2080
    id[food_apple_2081]=2081
    id[food_bacon_2082]=2082
    id[food_banana_2083]=2083
    id[food_bread_2084]=2084
    id[food_cake_2085]=2085
    id[food_carrot_2086]=2086
    id[food_cereal_2087]=2087
    id[food_cheese_2088]=2088
    id[food_chicken_2089]=2089
    id[food_dessert_2090]=2090
    id[food_donut_2091]=2091
    id[food_egg_2092]=2092
    id[food_fish_2093]=2093
    id[food_food_2094]=2094
    id[food_fruit_2095]=2095
    id[food_hamburger_2096]=2096
    id[food_ice_cream_2097]=2097
    id[food_jam_2098]=2098
    id[food_kiwi_2099]=2099
    id[food_lemon_2100]=2100
    id[food_noodles_2101]=2101
    id[food_oatmeal_2102]=2102
    id[food_orange_2103]=2103
    id[food_onion_2104]=2104
    id[food_peanut_butter_2105]=2105
    id[food_pizza_2106]=2106
    id[food_potato_2107]=2107
    id[food_rice_2108]=2108
    id[food_salt_2109]=2109
    id[food_snack_2110]=2110
    id[food_sugar_2111]=2111
    id[food_turkey_2112]=2112
    id[food_vegetable_2113]=2113
    id[dry_pasta_2114]=2114
    id[milk_2115]=2115
    id[clothes_dress_2116]=2116
    id[clothes_hat_2117]=2117
    id[clothes_gloves_2118]=2118
    id[clothes_jacket_2119]=2119
    id[clothes_scarf_2120]=2120
    id[clothes_underwear_2121]=2121
    id[knife_2122]=2122
    id[cutting_board_2123]=2123
    id[remote_control_2124]=2124
    id[soap_2125]=2125
    id[soap_2126]=2126
    id[towel_2128]=2128
    id[cd_player_2129]=2129
    id[dvd_player_2130]=2130
    id[headset_2131]=2131
    id[cup_2132]=2132
    id[cup_2133]=2133
    id[cup_2134]=2134
    id[stove_2135]=2135
    id[book_2136]=2136
    id[book_2137]=2137
    id[pot_2138]=2138
    id[vacuum_cleaner_2139]=2139
    id[bowl_2140]=2140
    id[bowl_2141]=2141
    id[bowl_2142]=2142
    id[cleaning_solution_2143]=2143
    id[ironing_board_2144]=2144
    id[cd_2145]=2145
    id[headset_2146]=2146
    id[phone_2147]=2147
    id[sauce_2148]=2148
    id[oil_2149]=2149
    id[fork_2150]=2150
    id[fork_2151]=2151
    id[plate_2152]=2152
    id[spectacles_2153]=2153
    id[fryingpan_2154]=2154
    id[detergent_2155]=2155
    id[window_2156]=2156
    id[bathroom_1]=1
    id[wall_2]=2
    id[wall_3]=3
    id[wall_4]=4
    id[wall_5]=5
    id[ceiling_6]=6
    id[ceiling_7]=7
    id[ceiling_8]=8
    id[ceiling_9]=9
    id[floor_10]=10
    id[floor_11]=11
    id[floor_12]=12
    id[floor_13]=13
    id[floor_14]=14
    id[toilet_15]=15
    id[shower_16]=16
    id[bathroom_cabinet_17]=17
    id[bathroom_counter_18]=18
    id[sink_19]=19
    id[faucet_20]=20
    id[shower_21]=21
    id[curtain_22]=22
    id[mat_32]=32
    id[drawing_33]=33
    id[walllamp_34]=34
    id[ceilinglamp_35]=35
    id[walllamp_36]=36
    id[doorjamb_37]=37
    id[door_38]=38
    id[light_39]=39
    id[dining_room_41]=41
    id[floor_42]=42
    id[floor_43]=43
    id[floor_44]=44
    id[floor_45]=45
    id[floor_46]=46
    id[floor_47]=47
    id[floor_48]=48
    id[floor_49]=49
    id[floor_50]=50
    id[floor_51]=51
    id[ceiling_52]=52
    id[ceiling_53]=53
    id[ceiling_54]=54
    id[ceiling_55]=55
    id[ceiling_56]=56
    id[ceiling_57]=57
    id[ceiling_58]=58
    id[ceiling_59]=59
    id[ceiling_60]=60
    id[door_61]=61
    id[door_62]=62
    id[wall_63]=63
    id[wall_64]=64
    id[wall_65]=65
    id[wall_66]=66
    id[wall_67]=67
    id[wall_68]=68
    id[wall_69]=69
    id[wall_70]=70
    id[phone_71]=71
    id[powersocket_72]=72
    id[light_73]=73
    id[knifeblock_76]=76
    id[pot_78]=78
    id[trashcan_99]=99
    id[mat_102]=102
    id[pillow_103]=103
    id[pillow_104]=104
    id[pillow_105]=105
    id[pillow_106]=106
    id[pillow_107]=107
    id[pillow_108]=108
    id[drawing_110]=110
    id[drawing_111]=111
    id[bench_113]=113
    id[table_114]=114
    id[bench_115]=115
    id[tvstand_116]=116
    id[cupboard_117]=117
    id[cupboard_118]=118
    id[kitchen_counter_119]=119
    id[sink_120]=120
    id[faucet_121]=121
    id[kitchen_counter_122]=122
    id[kitchen_counter_123]=123
    id[bookshelf_124]=124
    id[stovefan_125]=125
    id[fridge_126]=126
    id[oven_127]=127
    id[tray_128]=128
    id[dishwasher_129]=129
    id[coffe_maker_130]=130
    id[toaster_132]=132
    id[microwave_135]=135
    id[ceilinglamp_137]=137
    id[ceilinglamp_138]=138
    id[walllamp_139]=139
    id[walllamp_140]=140
    id[walllamp_141]=141
    id[bedroom_162]=162
    id[floor_163]=163
    id[floor_164]=164
    id[floor_165]=165
    id[floor_166]=166
    id[floor_167]=167
    id[floor_168]=168
    id[floor_169]=169
    id[floor_170]=170
    id[floor_171]=171
    id[floor_172]=172
    id[wall_173]=173
    id[wall_174]=174
    id[wall_175]=175
    id[wall_176]=176
    id[wall_177]=177
    id[wall_178]=178
    id[wall_179]=179
    id[wall_180]=180
    id[ceiling_181]=181
    id[ceiling_182]=182
    id[ceiling_183]=183
    id[ceiling_184]=184
    id[ceiling_185]=185
    id[ceiling_186]=186
    id[ceiling_187]=187
    id[ceiling_188]=188
    id[ceiling_189]=189
    id[doorjamb_190]=190
    id[window_191]=191
    id[nightstand_192]=192
    id[desk_193]=193
    id[chair_194]=194
    id[nightstand_195]=195
    id[bookshelf_196]=196
    id[bed_197]=197
    id[couch_198]=198
    id[table_199]=199
    id[filing_cabinet_200]=200
    id[drawing_201]=201
    id[drawing_202]=202
    id[mat_203]=203
    id[curtain_204]=204
    id[curtain_205]=205
    id[curtain_206]=206
    id[pillow_207]=207
    id[pillow_208]=208
    id[computer_209]=209
    id[cpuscreen_210]=210
    id[keyboard_211]=211
    id[light_212]=212
    id[mouse_213]=213
    id[mousepad_214]=214
    id[photoframe_219]=219
    id[ceilinglamp_237]=237
    id[tablelamp_238]=238
    id[tablelamp_239]=239
    id[home_office_241]=241
    id[wall_242]=242
    id[wall_243]=243
    id[wall_244]=244
    id[wall_245]=245
    id[wall_246]=246
    id[wall_247]=247
    id[wall_248]=248
    id[wall_249]=249
    id[ceiling_250]=250
    id[ceiling_251]=251
    id[ceiling_252]=252
    id[ceiling_253]=253
    id[ceiling_254]=254
    id[ceiling_255]=255
    id[ceiling_256]=256
    id[ceiling_257]=257
    id[ceiling_258]=258
    id[floor_259]=259
    id[floor_260]=260
    id[floor_261]=261
    id[floor_262]=262
    id[floor_263]=263
    id[floor_264]=264
    id[floor_265]=265
    id[floor_266]=266
    id[floor_267]=267
    id[floor_268]=268
    id[couch_269]=269
    id[table_270]=270
    id[chair_271]=271
    id[desk_272]=272
    id[tvstand_273]=273
    id[dresser_274]=274
    id[bookshelf_275]=275
    id[computer_276]=276
    id[cpuscreen_277]=277
    id[keyboard_278]=278
    id[mousepad_279]=279
    id[mouse_280]=280
    id[television_281]=281
    id[powersocket_282]=282
    id[light_283]=283
    id[mat_284]=284
    id[orchid_285]=285
    id[pillow_286]=286
    id[pillow_287]=287
    id[drawing_288]=288
    id[curtain_289]=289
    id[curtain_290]=290
    id[curtain_291]=291
    id[hanger_292]=292
    id[hanger_293]=293
    id[hanger_294]=294
    id[ceilinglamp_303]=303
    id[walllamp_304]=304
    id[walllamp_305]=305
    id[walllamp_306]=306
    id[walllamp_307]=307
    id[doorjamb_308]=308
    id[doorjamb_309]=309
    id[window_310]=310
    id[food_food_1000]=1000
    id[wooden_spoon_2000]=2000
    id[food_food_2001]=2001
    id[brush_2002]=2002
    id[chair_2003]=2003
    id[lighter_2004]=2004
    id[table_cloth_2005]=2005
    id[piano_bench_2006]=2006
    id[food_butter_2007]=2007
    id[diary_2008]=2008
    id[food_onion_2009]=2009
    id[soap_2010]=2010
    id[detergent_2011]=2011
    id[measuring_cup_2012]=2012
    id[oil_2013]=2013
    id[pencil_2014]=2014
    id[food_carrot_2015]=2015
    id[phone_2016]=2016
    id[phone_2017]=2017
    id[envelope_2018]=2018
    id[shampoo_2019]=2019
    id[pencil_2020]=2020
    id[food_food_2021]=2021
    id[stamp_2022]=2022
    id[tea_bag_2023]=2023
    id[ice_2024]=2024
    id[rag_2025]=2025
    id[check_2026]=2026
    id[food_orange_2027]=2027
    id[instrument_guitar_2028]=2028
    id[phone_2029]=2029
    id[cd_2030]=2030
    id[scrabble_2031]=2031
    id[shoes_2033]=2033
    id[laser_pointer_2034]=2034
    id[knife_2035]=2035
    id[clothes_pants_2036]=2036
    id[knife_2037]=2037
    id[box_2038]=2038
    id[lighter_2039]=2039
    id[pot_2040]=2040
    id[food_salt_2041]=2041
    id[after_shave_2042]=2042
    id[stamp_2043]=2043
    id[shoe_rack_2044]=2044
    id[glue_2045]=2045
    id[food_food_2046]=2046
    id[homework_2047]=2047
    id[food_onion_2048]=2048
    id[cup_2049]=2049
    id[stereo_2050]=2050
    id[after_shave_2051]=2051
    id[rag_2052]=2052
    id[coffee_filter_2053]=2053
    id[food_kiwi_2054]=2054
    id[envelope_2055]=2055
    id[toy_2056]=2056
    id[blow_dryer_2057]=2057
    id[check_2058]=2058
    id[tooth_paste_2059]=2059
    id[novel_2060]=2060
    id[food_orange_2061]=2061
    id[piano_bench_2062]=2062
    id[after_shave_2063]=2063
    id[food_food_2064]=2064
    id[coffee_filter_2065]=2065
    id[tea_2066]=2066
    id[piano_bench_2067]=2067
    id[tray_2068]=2068
    id[cat_2069]=2069
    id[chessboard_2070]=2070
    id[check_2071]=2071
    id[food_cheese_2072]=2072
    id[food_food_2073]=2073
    id[food_food_2074]=2074
    id[check_2075]=2075
    id[toilet_paper_2076]=2076
    id[food_peanut_butter_2077]=2077
    #id_end

    #size
    #size_end
