domain "virtualhome_debug"

typedef item: object
typedef character: object


#state
feature is_on(x: item)
feature is_off(x: item)
feature plugged(x: item)
feature unplugged(x: item)
feature open(x: item)
feature closed(x: item)
feature dirty(x: item)
feature clean(x: item)
feature sitting(x: character)
feature lying(x: character)

#add state
feature is_door(x: item)
feature is_explored(x: item)
feature is_room(x: item)

#relationship
feature on(x: item, y: item)
feature on_char(x: character, y: item)
feature inside(x: item, y: item)
feature inside_char(x: character, y: item)

feature between(x: item, y: item, z: item)
feature close_item(x: item, y: item)
feature close(x: character, y: item)
feature facing_item(x: item, y: item)
feature facing(x: character, y: item)
feature holds_rh(x: character, y: item)
feature holds_lh(x: character, y: item)

#Properties 
feature surfaces(x: item)
feature grabbable(x: item)
feature sittable(x: item)
feature lieable(x: item)
feature hangable(x: item)
feature drinkable(x: item)
feature eatable(x: item)
feature recipient(x: item)
feature cuttable(x: item)
feature pourable(x: item)
feature can_open(x: item)
feature has_switch(x: item)
feature readable(x: item)
feature lookable(x: item)
feature containers(x: item)
feature clothes(x: item)
feature person(x: item)
feature body_part(x: item)
feature cover_object(x: item)
feature has_plug(x: item)
feature has_paper(x: item)
feature movable(x: item)
feature cream(x: item)


object_constant char:character

#controllers
controller switchoff_executor(x: item)
controller switchon_executor(x: item)
controller put_executor(x: item, y: item)
controller grab_executor(x: item)
controller standup_executor(x: character)
controller wash_executor(x: item)
controller sit_executor(x: character)
controller open_executor(x: item)
controller close_executor(x: item)
controller pour_executor(x: item, y: item)
controller plugin_executor(x: item)
controller plugout_executor(x: item)
controller walk_executor(x: item)


def obj_inside_or_on(obj1: item, obj2: item):
  return inside(obj1, obj2) or on(obj2, obj1)

behavior walk(obj: item):
  goal: close(char, obj)
  body:
    walk_executor(obj)
  eff:
    foreach icf:item:
      if obj_inside_or_on(obj, icf):
        close[char, icf] = True