domain "virtualhome"

typedef item: object
typedef character: object

#  without return type annotations are assumed to be returning boolean values.

#state
on
off
plugged
unplugged
open
closed
dirty
clean
sitting(x: character)
lying(x: character)

#add state
room
comb
pillow
teeth
face_soap
sheets
mail
remote_control
instrument_violin
shoe_rack
lighter
food_vegetable
phone
table_cloth
pajamas
clothes_socks
form
face
wall_clock
food_egg
printing_paper
paper_towel
legs_both
glue
towel
coffee_table
food_sugar
microphone
foundation
curtain
mouse
duster
food_turkey
bookshelf
clothes_pants
food_onion
table
scrabble
wallshelf
sink
instrument_piano
food_snack
coin
tape
thread
towel_rack
electrical_outlet
dog
bathroom
hair
oil
sponge
cd_player
measuring_cup
food_apple
knifeblock
tablelamp
basket_for_clothes
drinking_glass
beer
novel
light_bulb
bathroom_cabinet
bench
dirt
food_orange
clothes_jacket
electric_shaver
envelope
coffee_cup
cleaning_solution
tea_bag
dough
longboard
napkin
clothes_skirt
walllamp
chef_knife
video_game_controller
detergent
hairdryer
balanceball
mirror
bedroom
mop
iron
shoes
cards
bag
fly
toilet
rag
clothes_shirt
fork
woman
closetdrawer
laser_pointer
deck_of_cards
food_noodles
razor
hands_both
drack
cup
console
food_cheese
video_game_console
bathroom_counter
kitchen_counter
oven
filing_cabinet
plate
brush
toaster
tooth_paste
shoe_shine_kit
pasta
toothbrush
keys
shelf
box
standingmirror
scors
board_game
mop_bucket
love_seat
bed
cloth_napkin
sauce_pan
drying_rack
ceilingfan
window
photoframe
facial_cleanser
cd
ceiling
dining_room
alarm_clock
floor_lamp
blender
stovefan
maindoor
band_aids
broom
food_dessert
food_bacon
check
diary
kettle
food_cake
ceilinglamp
bowl
spoon
chair
clothes_dress
dry_pasta
pantry
button
needle
food_donut
coffee_filter
piano_bench
microwave
food_bread
door
newspaper
food_salt
toilet_paper
coffee_pot
ground_coffee
food_pizza
headset
food_peanut_butter
man
food_ice_cream
laundry_detergent
cpuscreen
homework
bookmark
clothes_gloves
toothbrush_holder
ice
doorjamb
nightstand
alcohol
kitchen_cabinet
food_f
food_steak
dustpan
colander
washing_machine
food_jam
address_book
tvstand
dresser
candle
hanger
milk
food_carrot
cupboard
bathtub
purse
fax_machine
cleaning_bottle
tray
garbage_can
coffe_maker
instrument_guitar
food_food
floor
stamp
crayon
mousepad
oven_mitts
home_office
jelly
food_chicken
nail_pol
trashcan
clothes_scarf
cat
ironing_board
powersocket
televon
desk
food_cereal
spectacles
wine_glass
faucet
vacuum_cleaner
chessboard
child
food_oatmeal
d_soap
wooden_spoon
shampoo
dvd_player
music_stand
creditcard
centerpiece
food_rice
wine
couch
computer
orchid
stereo
vase
shredder
food_butter
mouthwash
after_shave
clothes_underwear
toy
knife
pot
keyboard
freezer
coffee
water_glass
drawing
shaving_cream
blow_dryer
soap
shower
picture
clothes_hat
wall
cutting_board
laptop
arms_both
pencil
dwasher
food_kiwi
water
conditioner
tea
hairbrush
feet_both
mat
juice
light
folder
bills


#relationship
on(x: item, y: item)
on_char(x: character, y: item)
inside(x: item, y: item)
inside_char(x: character, y: item)
between(door: item, room: item)
close(x: item, y: item)
close_char(x: character, y: item)
facing(x: item, y: item)
facing_char(x: character, y: item)
holds_rh(x: character, y: item)
holds_lh(x: character, y: item)

#Properties 
surfaces
grabbable
sittable
lieable
hangable
drinkable
eatable
recipient
cuttable
pourable
can_open
has_switch
readable
lookable
containers
clothes
person
body_part
cover_object
has_plug
has_paper
movable
cream


object_constant char:character

#
walk_executor
switchoff_executor
switchon_executor
put_executor(x: item, y: item)
grab_executor
standup_executor(x: character)
wash_executor
sit_executor(x: character)
open_executor
close_executor
pour_executor(x: item, y: item)
plugin_executor
plugout_executor


def inhand(inhand_obj:item):
  return holds_rh(char, inhand_obj) or holds_lh(char, inhand_obj)

def standing(char: character):
  return not sitting(char) and not lying(char)

def has_a_free_hand():
  symbol l=exs item1: item : holds_lh(char, item1)
  symbol r=exs item2: item : holds_rh(char, item2)
  return not l or not r



behavior put(inhand_obj: item, obj: item):
  body:
    assert surfaces(obj) or room(obj) or recipient(obj) or containers(obj) or can_open(obj)
    achieve inhand(inhand_obj)
    achieve close_char(char, obj)
    if can_open(obj) and closed(obj):
      achieve open(obj)
    put_executor(inhand_obj, obj)

  eff:
    holds_rh[char, inhand_obj] = False
    holds_lh[char, inhand_obj] = False
    if surfaces(obj):
      on[inhand_obj, obj] = True
    if room(obj) or recipient(obj) or containers(obj) or can_open(obj):
      inside[inhand_obj, obj] = True
    close[inhand_obj, obj] = True
    close[obj, inhand_obj] = True
    foreach inter:item:
      if close(inter, obj):
        close[inter, inhand_obj] = True
        close[inhand_obj, inter] = True
    if can_open(obj):
      open[obj] = True
      closed[obj] = False

behavior empty_a_hand():
  goal: has_a_free_hand()
  body:
    assert not has_a_free_hand()
    bind surf:item where:
      surfaces(surf)
    bind give_up_obj:item where:
      inhand(give_up_obj)
    put(give_up_obj, surf)

behavior stand():
  goal: standing(char)
  body:
    assert sitting(char) or lying(char)
    standup_executor(char)
  eff:
    sitting[char] = False
    lying[char] = False

behavior sit(obj: item):
  goal: sitting(char)
  body:
    assert not sitting(char)
    bind seat:item where:
      sittable(seat)
    achieve close_char(char, seat)
    sit_executor(seat)
  eff:
    sitting[char] = True
    on_char[char, seat] = True

def obj_inside_or_on(obj1: item, obj2: item):
  return inside(obj1, obj2) or on(obj2, obj1)

behavior walk(obj: item):
  goal: close_char(char, obj)
  body:
    achieve standing(char)
    walk_executor(obj)
  eff:
    foreach icf:item:
      close_char[char, icf]= False
      facing_char[char, icf]= False
      inside_char[char,icf]= False
      if obj_inside_or_on(obj, icf):
        close_char[char, icf] = True
    close_char[char,obj] = True

behavior switch_off(obj: item):
  goal: off(obj)
  body:
    assert has_switch(obj)
    assert on(obj)
    achieve has_a_free_hand()
    achieve close_char(char, obj)
    switchoff_executor(obj)
  eff:
    off[obj] = True
    on[obj] = False

behavior switch_on(obj: item):
  goal: on(obj)
  body:
    assert has_switch(obj)
    assert off(obj)
    achieve has_a_free_hand()
    achieve close_char(char, obj)
    switchon_executor(obj)
  eff:
    off[obj] = False
    on[obj] = True

behavior put_close(inhand_obj: item, obj: item):
  goal: close(inhand_obj, obj)
  body:
    put(inhand_obj, obj)

behavior put_on(inhand_obj: item, obj: item):
  goal: on(inhand_obj, obj)
  body:
    put(inhand_obj, obj)


behavior put_inside(inhand_obj: item, obj: item):
  goal: inside(inhand_obj, obj)
  body:
    put(inhand_obj, obj)

behavior grab(obj: item):
  goal: inhand(obj)
  body:
    assert grabbable(obj)
    achieve has_a_free_hand()
    foreach obj2:item:
      if inside(obj,obj2):
        if not room(obj2):
          assert can_open(obj2) or recipient(obj2)
          if can_open(obj2):
            achieve open(obj2)
    achieve close_char(char, obj)
    grab_executor(obj)
  eff:
    if exs item1: item : holds_lh(char, item1):
      holds_rh[char, obj] = True
    else:
      holds_lh[char, obj] = True

behavior wash(obj: item):
  goal: clean(obj)
  body:
    achieve has_a_free_hand()
    achieve close_char(char, obj)
    wash_executor(obj)
  eff:
    dirty[obj] = False
    clean[obj] = True

behavior open(obj: item):
  goal: open(obj)
  body:
    assert can_open(obj)
    assert closed(obj)
    achieve has_a_free_hand()
    achieve close_char(char, obj)
    open_executor(obj)
  eff:
    open[obj] = True
    closed[obj] = False

behavior close(obj: item):
  goal: closed(obj)
  body:
    assert can_open(obj)
    assert open(obj)
    achieve has_a_free_hand()
    achieve close_char(char, obj)
    close_executor(obj)
  eff:
    open[obj] = False
    closed[obj] = True

behavior pour(obj: item, target: item):
  goal: inside(obj, target)
  body:
    assert pourable(obj) or drinkable(obj)
    assert recipient(target)
    achieve inhand(obj)
    achieve close_char(char, target)
    pour_executor(obj, target)
  eff:
    inside[obj, target] = True

behavior plugin(object:item):
  goal: plugged(object)
  body:
    assert has_plug(object)
    assert unplugged(object)
    achieve has_a_free_hand()
    achieve close_char(char, object)
    plugin_executor(object)
  eff:
    plugged[object] = True
    unplugged[object] = False
  
behavior plugout(object:item):
  goal: unplugged(object)
  body:
    assert has_plug(object)
    assert plugged(object)
    achieve has_a_free_hand()
    achieve close_char(char, object)
    plugout_executor(object)
  eff:
    plugged[object] = False
    unplugged[object] = True