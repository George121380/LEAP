Make Chicken Stir-Fry.
Cut chicken into thin strips and season with salt and pepper.In a pan, heat oil over. Add minced garlic and ginger, then the chicken. Add mixed vegetables and stir-fry until tender-crisp.

behavior prepare_chicken(chicken:item, salt:item, pepper:item):
    body:
        achieve sliced(chicken)
        achieve inside(salt, chicken)
        achieve inside(pepper, chicken)

behavior start_stove(stove:item):
    body:
        achieve is_on(stove)

behavior heat_oil_on_pan(pan:item, stove:item, oil:item):
    body:
        achieve on(pan, stove)
        start_stove(stove)
        achieve inside(oil, pan)

behavior cook_chicken_with_garlic_ginger(pan:item, chicken:item, garlic:item, ginger:item):
    body:
        achieve inside(garlic, pan)
        achieve inside(ginger, pan)
        achieve inside(chicken, pan)
        achieve fried(chicken)

behavior add_vegetables_and_stir_fry(pan:item, stove:item, vegetables:item):
    body:
        achieve inside(vegetables, pan)
        achieve is_on(stove)

behavior __goal__():
    body:
        bind stove: item where:
            is_stove(stove)
        bind pan: item where:
            is_pan(pan)
        bind chicken: item where:
            is_chicken(chicken)
        bind oil: item where:
            is_oil(oil)
        bind salt: item where:
            is_salt(salt)
        bind pepper: item where:
            is_pepper(pepper)
        bind garlic: item where:
            is_garlic(garlic)
        bind ginger: item where:
            is_ginger(ginger)
        bind vegetables: item where:
            is_tomato(vegetables)
        prepare_chicken(chicken, salt, pepper)
        heat_oil_on_pan(pan, stove, oil)
        cook_chicken_with_garlic_ginger(pan, chicken, garlic, ginger)
        add_vegetables_and_stir_fry(pan, stove, vegetables)