problem "agent-problem"
domain "kitchen_partial_ability.cdl"

#!pragma planner_is_goal_serializable=False
#!pragma planner_is_goal_ordered=True
#!pragma planner_always_commit_skeleton=True

objects:
  tomato_1:item
  tomato_2:item
  tomato_3:item
  tomato_4:item
  egg_5:item
  egg_6:item
  egg_7:item
  egg_8:item
  oil_9:item
  sugar_10:item
  pan_11:item
  salt_12:item
  bowl_13:item
  bowl_14:item
  bowl_15:item
  bowl_16:item
  knife_17:item
  fridge_18:item
  stove_19:item
  sink_20:item
  faucet_21:item
  spatula_22:item
  countertop_23:item
  water_24:item
  pepper_25:item
  bread_26:item
  onion_27:item
  bacon_28:item
  cheese_29:item
  bread_30:item
  bread_31:item
  bread_32:item
  pot_33:item
  noodles_34:item
  chicken_35:item
  garlic_36:item
  ginger_37:item
  vegetables_38:item
  oven_39:item
  plate_40:item
  plate_41:item
  plate_42:item
  plate_43:item
  cuttingboard_44:item
  beef_45:item
  potato_46:item
  shrimp_47:item
#object_end

init:
    #categories
    is_tomato[tomato_1]=True
    is_tomato[tomato_2]=True
    is_tomato[tomato_3]=True
    is_tomato[tomato_4]=True
    is_egg[egg_5]=True
    is_egg[egg_6]=True
    is_egg[egg_7]=True
    is_egg[egg_8]=True
    is_oil[oil_9]=True
    is_sugar[sugar_10]=True
    is_pan[pan_11]=True
    is_salt[salt_12]=True
    is_bowl[bowl_13]=True
    is_bowl[bowl_14]=True
    is_bowl[bowl_15]=True
    is_bowl[bowl_16]=True
    is_knife[knife_17]=True
    is_fridge[fridge_18]=True
    is_stove[stove_19]=True
    is_sink[sink_20]=True
    is_faucet[faucet_21]=True
    is_spatula[spatula_22]=True
    is_countertop[countertop_23]=True
    is_water[water_24]=True
    is_pepper[pepper_25]=True
    is_bread[bread_26]=True
    is_onion[onion_27]=True
    is_bacon[bacon_28]=True
    is_cheese[cheese_29]=True
    is_bread[bread_30]=True
    is_bread[bread_31]=True
    is_bread[bread_32]=True
    is_pot[pot_33]=True
    is_noodles[noodles_34]=True
    is_chicken[chicken_35]=True
    is_garlic[garlic_36]=True
    is_ginger[ginger_37]=True
    is_vegetables[vegetables_38]=True
    is_oven[oven_39]=True
    is_plate[plate_40]=True
    is_plate[plate_41]=True
    is_plate[plate_42]=True
    is_plate[plate_43]=True
    is_cuttingboard[cuttingboard_44]=True
    is_beef[beef_45]=True
    is_potato[potato_46]=True
    is_shrimp[shrimp_47]=True
    #categories_end

    #states
    is_off[stove_19]=True
    is_off[faucet_21]=True
    is_off[oven_39]=True
    closed[fridge_18]=True
    closed[oven_39]=True
    dirty[tomato_1]=True
    dirty[tomato_2]=True
    dirty[tomato_3]=True
    dirty[tomato_4]=True
    dirty[onion_27]=True
    dirty[vegetables_38]=True
    clean[pan_11]=True
    clean[bowl_13]=True
    clean[bowl_14]=True
    clean[bowl_15]=True
    clean[bowl_16]=True
    clean[pot_33]=True
    clean[plate_40]=True
    clean[plate_41]=True
    clean[plate_42]=True
    clean[plate_43]=True
    #states_end

    #char
    #char_end

    #properties
    surfaces[stove_19]=True
    surfaces[countertop_23]=True
    surfaces[cuttingboard_44]=True
    grabbable[tomato_1]=True
    grabbable[tomato_2]=True
    grabbable[tomato_3]=True
    grabbable[tomato_4]=True
    grabbable[egg_5]=True
    grabbable[egg_6]=True
    grabbable[egg_7]=True
    grabbable[egg_8]=True
    grabbable[oil_9]=True
    grabbable[sugar_10]=True
    grabbable[pan_11]=True
    grabbable[salt_12]=True
    grabbable[bowl_13]=True
    grabbable[bowl_14]=True
    grabbable[bowl_15]=True
    grabbable[bowl_16]=True
    grabbable[knife_17]=True
    grabbable[spatula_22]=True
    grabbable[pepper_25]=True
    grabbable[bread_26]=True
    grabbable[onion_27]=True
    grabbable[bacon_28]=True
    grabbable[cheese_29]=True
    grabbable[bread_30]=True
    grabbable[bread_31]=True
    grabbable[bread_32]=True
    grabbable[pot_33]=True
    grabbable[noodles_34]=True
    grabbable[chicken_35]=True
    grabbable[garlic_36]=True
    grabbable[ginger_37]=True
    grabbable[vegetables_38]=True
    grabbable[plate_40]=True
    grabbable[plate_41]=True
    grabbable[plate_42]=True
    grabbable[plate_43]=True
    grabbable[cuttingboard_44]=True
    grabbable[beef_45]=True
    grabbable[potato_46]=True
    grabbable[shrimp_47]=True
    cuttable[tomato_1]=True
    cuttable[tomato_2]=True
    cuttable[tomato_3]=True
    cuttable[tomato_4]=True
    cuttable[bread_26]=True
    cuttable[onion_27]=True
    cuttable[bacon_28]=True
    cuttable[cheese_29]=True
    cuttable[bread_30]=True
    cuttable[bread_31]=True
    cuttable[bread_32]=True
    cuttable[noodles_34]=True
    cuttable[chicken_35]=True
    cuttable[garlic_36]=True
    cuttable[ginger_37]=True
    cuttable[vegetables_38]=True
    cuttable[beef_45]=True
    cuttable[potato_46]=True
    cuttable[shrimp_47]=True
    pourable[salt_12]=True
    pourable[pepper_25]=True
    can_open[fridge_18]=True
    can_open[oven_39]=True
    has_switch[stove_19]=True
    has_switch[faucet_21]=True
    has_switch[oven_39]=True
    containers[pan_11]=True
    containers[bowl_13]=True
    containers[bowl_14]=True
    containers[bowl_15]=True
    containers[bowl_16]=True
    containers[fridge_18]=True
    containers[sink_20]=True
    containers[pot_33]=True
    containers[oven_39]=True
    containers[plate_40]=True
    containers[plate_41]=True
    containers[plate_42]=True
    containers[plate_43]=True
    peelable[tomato_1]=True
    peelable[tomato_2]=True
    peelable[tomato_3]=True
    peelable[tomato_4]=True
    peelable[potato_46]=True
    peelable[shrimp_47]=True
    storable[countertop_23]=True
    eatable[tomato_1]=True
    eatable[tomato_2]=True
    eatable[tomato_3]=True
    eatable[tomato_4]=True
    eatable[egg_5]=True
    eatable[egg_6]=True
    eatable[egg_7]=True
    eatable[egg_8]=True
    eatable[oil_9]=True
    eatable[sugar_10]=True
    eatable[salt_12]=True
    eatable[pepper_25]=True
    eatable[bread_26]=True
    eatable[onion_27]=True
    eatable[bacon_28]=True
    eatable[cheese_29]=True
    eatable[bread_30]=True
    eatable[bread_31]=True
    eatable[bread_32]=True
    eatable[noodles_34]=True
    eatable[chicken_35]=True
    eatable[garlic_36]=True
    eatable[ginger_37]=True
    eatable[vegetables_38]=True
    eatable[beef_45]=True
    eatable[potato_46]=True
    eatable[shrimp_47]=True
    cookaware[pan_11]=True
    cookaware[pot_33]=True
    cookaware[oven_39]=True
    #properties_end

    #relations
    on[faucet_21,sink_20]=True
    on[oven_39,countertop_23]=True
    close[sink_20,faucet_21]=True
    close[faucet_21,sink_20]=True
    close[countertop_23,oven_39]=True
    close[oven_39,countertop_23]=True
    #relations_end

    #exploration
    known[fridge_18]=True
    known[stove_19]=True
    known[sink_20]=True
    known[faucet_21]=True
    known[countertop_23]=True
    known[oven_39]=True
    #exploration_end

    #id
    id[tomato_1]=1
    id[tomato_2]=2
    id[tomato_3]=3
    id[tomato_4]=4
    id[egg_5]=5
    id[egg_6]=6
    id[egg_7]=7
    id[egg_8]=8
    id[oil_9]=9
    id[sugar_10]=10
    id[pan_11]=11
    id[salt_12]=12
    id[bowl_13]=13
    id[bowl_14]=14
    id[bowl_15]=15
    id[bowl_16]=16
    id[knife_17]=17
    id[fridge_18]=18
    id[stove_19]=19
    id[sink_20]=20
    id[faucet_21]=21
    id[spatula_22]=22
    id[countertop_23]=23
    id[water_24]=24
    id[pepper_25]=25
    id[bread_26]=26
    id[onion_27]=27
    id[bacon_28]=28
    id[cheese_29]=29
    id[bread_30]=30
    id[bread_31]=31
    id[bread_32]=32
    id[pot_33]=33
    id[noodles_34]=34
    id[chicken_35]=35
    id[garlic_36]=36
    id[ginger_37]=37
    id[vegetables_38]=38
    id[oven_39]=39
    id[plate_40]=40
    id[plate_41]=41
    id[plate_42]=42
    id[plate_43]=43
    id[cuttingboard_44]=44
    id[beef_45]=45
    id[potato_46]=46
    id[shrimp_47]=47
    #id_end

#goal_representation
## Series of formal representations of find actions

behavior find_onion_27_in_countertop_23(onion27:item):
    goal: known(onion27)
    body:
        assert is_onion(onion27)
        bind countertop23:item where:
            is_countertop(countertop23) and id(countertop23)==23
        achieve close_char(char,countertop23)
    eff:
        foreach o:item:
            if is_onion(o):
                known[o] = True
                on[o,countertop23] = True

behavior find_potato_46_in_countertop_23(potato46:item):
    goal: known(potato46)
    body:
        assert is_potato(potato46)
        bind countertop23:item where:
            is_countertop(countertop23) and id(countertop23)==23
        achieve close_char(char,countertop23)
    eff:
        foreach o:item:
            if is_potato(o):
                known[o] = True
                on[o,countertop23] = True

behavior find_bread_31_in_countertop_23(bread31:item):
    goal: known(bread31)
    body:
        assert is_bread(bread31)
        bind countertop23:item where:
            is_countertop(countertop23) and id(countertop23)==23
        achieve close_char(char,countertop23)
    eff:
        foreach o:item:
            if is_bread(o):
                known[o] = True
                on[o,countertop23] = True

behavior find_bacon_28_in_fridge_18(bacon28:item):
    goal: known(bacon28)
    body:
        assert is_bacon(bacon28)
        bind fridge18:item where:
            is_fridge(fridge18) and id(fridge18)==18
        achieve close_char(char,fridge18)
        achieve open(fridge18)
    eff:
        foreach o:item:
            if is_bacon(o):
                known[o] = True
                inside[o,fridge18] = True
                
behavior find_oil_9_in_countertop_23(oil9:item):
    goal: known(oil9)
    body:
        assert is_oil(oil9)
        bind countertop23:item where:
            is_countertop(countertop23) and id(countertop23)==23
        achieve close_char(char,countertop23)
    eff:
        foreach o:item:
            if is_oil(o):
                known[o] = True
                on[o,countertop23] = True

behavior find_ginger_37_in_countertop_23(ginger37:item):
    goal: known(ginger37)
    body:
        assert is_ginger(ginger37)
        bind countertop23:item where:
            is_countertop(countertop23) and id(countertop23)==23
        achieve close_char(char,countertop23)
    eff:
        foreach o:item:
            if is_ginger(o):
                known[o] = True
                on[o,countertop23] = True

behavior find_cheese_29_in_fridge_18(cheese29:item):
    goal: known(cheese29)
    body:
        assert is_cheese(cheese29)
        bind fridge18:item where:
            is_fridge(fridge18) and id(fridge18)==18
        achieve close_char(char,fridge18)
        achieve open(fridge18)
    eff:
        foreach o:item:
            if is_cheese(o):
                known[o] = True
                inside[o,fridge18] = True

behavior find_plate_43_in_countertop_23(plate43:item):
    goal: known(plate43)
    body:
        assert is_plate(plate43)
        bind countertop23:item where:
            is_countertop(countertop23) and id(countertop23)==23
        achieve close_char(char,countertop23)
    eff:
        foreach o:item:
            if is_plate(o):
                known[o] = True
                on[o,countertop23] = True
                
behavior find_bowl_16_in_countertop_23(bowl16:item):
    goal: known(bowl16)
    body:
        assert is_bowl(bowl16)
        bind countertop23:item where:
            is_countertop(countertop23) and id(countertop23)==23
        achieve close_char(char,countertop23)
    eff:
        foreach o:item:
            if is_bowl(o):
                known[o] = True
                on[o,countertop23] = True

behavior find_vegetables_38_in_fridge_18(vegetables38:item):
    goal: known(vegetables38)
    body:
        assert is_vegetables(vegetables38)
        bind fridge18:item where:
            is_fridge(fridge18) and id(fridge18)==18
        achieve close_char(char,fridge18)
        achieve open(fridge18)
    eff:
        foreach o:item:
            if is_vegetables(o):
                known[o] = True
                inside[o,fridge18] = True
                
behavior find_shrimp_47_in_fridge_18(shrimp47:item):
    goal: known(shrimp47)
    body:
        assert is_shrimp(shrimp47)
        bind fridge18:item where:
            is_fridge(fridge18) and id(fridge18)==18
        achieve close_char(char,fridge18)
        achieve open(fridge18)
    eff:
        foreach o:item:
            if is_shrimp(o):
                known[o] = True
                inside[o,fridge18] = True

behavior find_pan_11_in_stove_19(pan11:item):
    goal: known(pan11)
    body:
        assert is_pan(pan11)
        bind stove19:item where:
            is_stove(stove19) and id(stove19) == 19
        achieve close_char(char,stove19)
    eff:
        foreach o:item:
            if is_pan(o):
                known[o] = True
                on[o,stove19] = True

behavior find_noodles_34_in_countertop_23(noodles34:item):
    goal: known(noodles34)
    body:
        assert is_noodles(noodles34)
        bind countertop23:item where:
            is_countertop(countertop23) and id(countertop23) == 23
        achieve close_char(char,countertop23)
    eff:
        foreach o:item:
            if is_noodles(o):
                known[o] = True
                on[o,countertop23] = True

behavior find_egg_7_in_fridge_18(egg7:item):
    goal: known(egg7)
    body:
        assert is_egg(egg7)
        bind fridge18:item where:
            is_fridge(fridge18) and id(fridge18) == 18
        achieve close_char(char,fridge18)
        achieve open(fridge18)
    eff:
        foreach o:item:
            if is_egg(o):
                known[o] = True
                inside[o,fridge18] = True

behavior find_spatula_22_in_countertop_23(spatula22:item):
    goal: known(spatula22)
    body:
        assert is_spatula(spatula22)
        bind countertop23:item where:
            is_countertop(countertop23) and id(countertop23) == 23
        achieve close_char(char,countertop23)
    eff:
        foreach o:item:
            if is_spatula(o):
                known[o] = True
                on[o,countertop23] = True

behavior find_beef_45_in_fridge_18(beef45:item):
    goal: known(beef45)
    body:
        assert is_beef(beef45)
        bind fridge18:item where:
            is_fridge(fridge18) and id(fridge18)==18
        achieve close_char(char,fridge18)
        achieve open(fridge18)
    eff:
        foreach o:item:
            if is_beef(o):
                known[o] = True
                inside[o,fridge18] = True

behavior find_pepper_25_in_countertop_23(pepper25:item):
    goal: known(pepper25)
    body:
        assert is_pepper(pepper25)
        bind countertop23:item where:
            is_countertop(countertop23) and id(countertop23) == 23
        achieve close_char(char,countertop23)
    eff:
        foreach o:item:
            if is_pepper(o):
                known[o] = True
                on[o,countertop23] = True

behavior find_pot_33_in_countertop_23(pot33:item):
    goal: known(pot33)
    body:
        assert is_pot(pot33)
        bind countertop23:item where:
            is_countertop(countertop23) and id(countertop23) == 23
        achieve close_char(char,countertop23)
    eff:
        foreach o:item:
            if is_pot(o):
                known[o] = True
                on[o,countertop23] = True

behavior find_chicken_35_in_fridge_18(chicken35:item):
    goal: known(chicken35)
    body:
        assert is_chicken(chicken35)
        bind fridge18:item where:
            is_fridge(fridge18) and id(fridge18)==18
        achieve close_char(char,fridge18)
        achieve open(fridge18)
    eff:
        foreach o:item:
            if is_chicken(o):
                known[o] = True
                inside[o,fridge18] = True

behavior find_cuttingboard_44_in_countertop_23(cuttingboard44:item):
    goal: known(cuttingboard44)
    body:
        assert is_cuttingboard(cuttingboard44)
        bind countertop23:item where:
            is_countertop(countertop23) and id(countertop23)==23
        achieve close_char(char,countertop23)
    eff:
        foreach o:item:
            if is_cuttingboard(o):
                known[o] = True
                on[o,countertop23] = True

behavior find_garlic_36_in_countertop_23(garlic36:item):
    goal: known(garlic36)
    body:
        assert is_garlic(garlic36)
        bind countertop23:item where:
            is_countertop(countertop23) and id(countertop23) == 23
        achieve close_char(char,countertop23)
    eff:
        foreach o:item:
            if is_garlic(o):
                known[o] = True
                on[o,countertop23] = True

behavior find_water_24_in_sink_20(water24:item):
    goal: known(water24)
    body:
        assert is_water(water24)
        bind sink20:item where:
            is_sink(sink20) and id(sink20)==20
        achieve close_char(char,sink20)
    eff:
        foreach o:item:
            if is_water(o):
                known[o] = True
                inside[o,sink20] = True

behavior find_knife_17_in_countertop_23(knife17:item):
    goal: known(knife17)
    body:
        assert is_knife(knife17) 
        bind countertop23:item where:
            is_countertop(countertop23) and id(countertop23)==23
        achieve close_char(char,countertop23)
    eff:
        foreach o:item:
            if is_knife(o):
                known[o] = True
                on[o,countertop23] = True

behavior find_sugar_10_in_countertop_23(sugar10:item):
    goal: known(sugar10)
    body:
        assert is_sugar(sugar10)
        bind countertop23:item where:
            is_countertop(countertop23) and id(countertop23) == 23
        achieve close_char(char,countertop23)
    eff:
        foreach o:item:
            if is_sugar(o):
                known[o] = True
                on[o,countertop23] = True

behavior find_tomato_1_in_countertop_23(tomato1:item):
    goal: known(tomato1)
    body:
        assert is_tomato(tomato1)
        bind countertop23:item where:
            is_countertop(countertop23) and id(countertop23) == 23
        achieve close_char(char,countertop23)
    eff:
        foreach o:item:
            if is_tomato(o):
                known[o] = True
                on[o,countertop23] = True

behavior find_salt_12_in_countertop_23(salt12:item):
    goal: known(salt12)
    body:
        assert is_salt(salt12)
        bind countertop23:item where:
            is_countertop(countertop23) and id(countertop23) == 23
        achieve close_char(char,countertop23)
    eff:
        foreach o:item:
            if is_salt(o):
                known[o] = True
                on[o,countertop23] = True

behavior clean_object(obj: item):
    goal: clean(obj)
    body:
        bind sink: item where:
            is_sink(sink)
        bind faucet: item where:
            is_faucet(faucet)
        achieve inside(obj, sink)
        achieve_once is_on(faucet)
        achieve clean(obj)
        achieve_once is_off(faucet)

behavior prepare_bacon_cheese_tomato_sandwich(bacon:item, cheese:item, tomato:item, sandwich:item):
    body:
        achieve clean(bacon)
        achieve clean(cheese)
        achieve clean(tomato)
        achieve sliced(tomato)
        achieve inside(bacon, sandwich)
        achieve inside(cheese, sandwich)
        achieve inside(tomato, sandwich)

behavior __goal__():
    body:
        bind bacon: item where:
            is_bacon(bacon)
        bind cheese: item where:
            is_cheese(cheese)
        bind tomato: item where:
            is_tomato(tomato)
        bind sandwich: item where:
            is_bread(sandwich)
        clean_object(bacon)
        clean_object(cheese)
        clean_object(tomato)
        prepare_bacon_cheese_tomato_sandwich(bacon, cheese, tomato, sandwich)

#goal_representation_end
