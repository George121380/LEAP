 
behavior find_pot(pot:item):
    body:
        achieve_once inhand(pot)

behavior fill_pot_with_water(pot:item):
    body:
        achieve has_water(pot)

behavior put_pot_on_stove(pot:item, stove:item):
    body:
        achieve on(pot, stove)

behavior __goal__():
    body:
        bind pot: item where:
            is_pot(pot)
        # Select a pot
        
        bind stove: item where:
            is_stove(stove)
        # Select a stove

        find_pot(pot)
        fill_pot_with_water(pot)
        put_pot_on_stove(pot, stove)
